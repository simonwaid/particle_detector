magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< error_p >>
rect -678 581 -620 587
rect -560 581 -502 587
rect -442 581 -384 587
rect -324 581 -266 587
rect -206 581 -148 587
rect -88 581 -30 587
rect 30 581 88 587
rect 148 581 206 587
rect 266 581 324 587
rect 384 581 442 587
rect 502 581 560 587
rect 620 581 678 587
rect -678 547 -666 581
rect -560 547 -548 581
rect -442 547 -430 581
rect -324 547 -312 581
rect -206 547 -194 581
rect -88 547 -76 581
rect 30 547 42 581
rect 148 547 160 581
rect 266 547 278 581
rect 384 547 396 581
rect 502 547 514 581
rect 620 547 632 581
rect -678 541 -620 547
rect -560 541 -502 547
rect -442 541 -384 547
rect -324 541 -266 547
rect -206 541 -148 547
rect -88 541 -30 547
rect 30 541 88 547
rect 148 541 206 547
rect 266 541 324 547
rect 384 541 442 547
rect 502 541 560 547
rect 620 541 678 547
rect -678 71 -620 77
rect -560 71 -502 77
rect -442 71 -384 77
rect -324 71 -266 77
rect -206 71 -148 77
rect -88 71 -30 77
rect 30 71 88 77
rect 148 71 206 77
rect 266 71 324 77
rect 384 71 442 77
rect 502 71 560 77
rect 620 71 678 77
rect -678 37 -666 71
rect -560 37 -548 71
rect -442 37 -430 71
rect -324 37 -312 71
rect -206 37 -194 71
rect -88 37 -76 71
rect 30 37 42 71
rect 148 37 160 71
rect 266 37 278 71
rect 384 37 396 71
rect 502 37 514 71
rect 620 37 632 71
rect -678 31 -620 37
rect -560 31 -502 37
rect -442 31 -384 37
rect -324 31 -266 37
rect -206 31 -148 37
rect -88 31 -30 37
rect 30 31 88 37
rect 148 31 206 37
rect 266 31 324 37
rect 384 31 442 37
rect 502 31 560 37
rect 620 31 678 37
rect -678 -37 -620 -31
rect -560 -37 -502 -31
rect -442 -37 -384 -31
rect -324 -37 -266 -31
rect -206 -37 -148 -31
rect -88 -37 -30 -31
rect 30 -37 88 -31
rect 148 -37 206 -31
rect 266 -37 324 -31
rect 384 -37 442 -31
rect 502 -37 560 -31
rect 620 -37 678 -31
rect -678 -71 -666 -37
rect -560 -71 -548 -37
rect -442 -71 -430 -37
rect -324 -71 -312 -37
rect -206 -71 -194 -37
rect -88 -71 -76 -37
rect 30 -71 42 -37
rect 148 -71 160 -37
rect 266 -71 278 -37
rect 384 -71 396 -37
rect 502 -71 514 -37
rect 620 -71 632 -37
rect -678 -77 -620 -71
rect -560 -77 -502 -71
rect -442 -77 -384 -71
rect -324 -77 -266 -71
rect -206 -77 -148 -71
rect -88 -77 -30 -71
rect 30 -77 88 -71
rect 148 -77 206 -71
rect 266 -77 324 -71
rect 384 -77 442 -71
rect 502 -77 560 -71
rect 620 -77 678 -71
rect -678 -547 -620 -541
rect -560 -547 -502 -541
rect -442 -547 -384 -541
rect -324 -547 -266 -541
rect -206 -547 -148 -541
rect -88 -547 -30 -541
rect 30 -547 88 -541
rect 148 -547 206 -541
rect 266 -547 324 -541
rect 384 -547 442 -541
rect 502 -547 560 -541
rect 620 -547 678 -541
rect -678 -581 -666 -547
rect -560 -581 -548 -547
rect -442 -581 -430 -547
rect -324 -581 -312 -547
rect -206 -581 -194 -547
rect -88 -581 -76 -547
rect 30 -581 42 -547
rect 148 -581 160 -547
rect 266 -581 278 -547
rect 384 -581 396 -547
rect 502 -581 514 -547
rect 620 -581 632 -547
rect -678 -587 -620 -581
rect -560 -587 -502 -581
rect -442 -587 -384 -581
rect -324 -587 -266 -581
rect -206 -587 -148 -581
rect -88 -587 -30 -581
rect 30 -587 88 -581
rect 148 -587 206 -581
rect 266 -587 324 -581
rect 384 -587 442 -581
rect 502 -587 560 -581
rect 620 -587 678 -581
<< pwell >>
rect -875 -719 875 719
<< nmoslvt >>
rect -679 109 -619 509
rect -561 109 -501 509
rect -443 109 -383 509
rect -325 109 -265 509
rect -207 109 -147 509
rect -89 109 -29 509
rect 29 109 89 509
rect 147 109 207 509
rect 265 109 325 509
rect 383 109 443 509
rect 501 109 561 509
rect 619 109 679 509
rect -679 -509 -619 -109
rect -561 -509 -501 -109
rect -443 -509 -383 -109
rect -325 -509 -265 -109
rect -207 -509 -147 -109
rect -89 -509 -29 -109
rect 29 -509 89 -109
rect 147 -509 207 -109
rect 265 -509 325 -109
rect 383 -509 443 -109
rect 501 -509 561 -109
rect 619 -509 679 -109
<< ndiff >>
rect -737 497 -679 509
rect -737 121 -725 497
rect -691 121 -679 497
rect -737 109 -679 121
rect -619 497 -561 509
rect -619 121 -607 497
rect -573 121 -561 497
rect -619 109 -561 121
rect -501 497 -443 509
rect -501 121 -489 497
rect -455 121 -443 497
rect -501 109 -443 121
rect -383 497 -325 509
rect -383 121 -371 497
rect -337 121 -325 497
rect -383 109 -325 121
rect -265 497 -207 509
rect -265 121 -253 497
rect -219 121 -207 497
rect -265 109 -207 121
rect -147 497 -89 509
rect -147 121 -135 497
rect -101 121 -89 497
rect -147 109 -89 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 89 497 147 509
rect 89 121 101 497
rect 135 121 147 497
rect 89 109 147 121
rect 207 497 265 509
rect 207 121 219 497
rect 253 121 265 497
rect 207 109 265 121
rect 325 497 383 509
rect 325 121 337 497
rect 371 121 383 497
rect 325 109 383 121
rect 443 497 501 509
rect 443 121 455 497
rect 489 121 501 497
rect 443 109 501 121
rect 561 497 619 509
rect 561 121 573 497
rect 607 121 619 497
rect 561 109 619 121
rect 679 497 737 509
rect 679 121 691 497
rect 725 121 737 497
rect 679 109 737 121
rect -737 -121 -679 -109
rect -737 -497 -725 -121
rect -691 -497 -679 -121
rect -737 -509 -679 -497
rect -619 -121 -561 -109
rect -619 -497 -607 -121
rect -573 -497 -561 -121
rect -619 -509 -561 -497
rect -501 -121 -443 -109
rect -501 -497 -489 -121
rect -455 -497 -443 -121
rect -501 -509 -443 -497
rect -383 -121 -325 -109
rect -383 -497 -371 -121
rect -337 -497 -325 -121
rect -383 -509 -325 -497
rect -265 -121 -207 -109
rect -265 -497 -253 -121
rect -219 -497 -207 -121
rect -265 -509 -207 -497
rect -147 -121 -89 -109
rect -147 -497 -135 -121
rect -101 -497 -89 -121
rect -147 -509 -89 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 89 -121 147 -109
rect 89 -497 101 -121
rect 135 -497 147 -121
rect 89 -509 147 -497
rect 207 -121 265 -109
rect 207 -497 219 -121
rect 253 -497 265 -121
rect 207 -509 265 -497
rect 325 -121 383 -109
rect 325 -497 337 -121
rect 371 -497 383 -121
rect 325 -509 383 -497
rect 443 -121 501 -109
rect 443 -497 455 -121
rect 489 -497 501 -121
rect 443 -509 501 -497
rect 561 -121 619 -109
rect 561 -497 573 -121
rect 607 -497 619 -121
rect 561 -509 619 -497
rect 679 -121 737 -109
rect 679 -497 691 -121
rect 725 -497 737 -121
rect 679 -509 737 -497
<< ndiffc >>
rect -725 121 -691 497
rect -607 121 -573 497
rect -489 121 -455 497
rect -371 121 -337 497
rect -253 121 -219 497
rect -135 121 -101 497
rect -17 121 17 497
rect 101 121 135 497
rect 219 121 253 497
rect 337 121 371 497
rect 455 121 489 497
rect 573 121 607 497
rect 691 121 725 497
rect -725 -497 -691 -121
rect -607 -497 -573 -121
rect -489 -497 -455 -121
rect -371 -497 -337 -121
rect -253 -497 -219 -121
rect -135 -497 -101 -121
rect -17 -497 17 -121
rect 101 -497 135 -121
rect 219 -497 253 -121
rect 337 -497 371 -121
rect 455 -497 489 -121
rect 573 -497 607 -121
rect 691 -497 725 -121
<< psubdiff >>
rect -839 649 -743 683
rect 743 649 839 683
rect -839 587 -805 649
rect 805 587 839 649
rect -839 -649 -805 -587
rect 805 -649 839 -587
rect -839 -683 -743 -649
rect 743 -683 839 -649
<< psubdiffcont >>
rect -743 649 743 683
rect -839 -587 -805 587
rect 805 -587 839 587
rect -743 -683 743 -649
<< poly >>
rect -682 581 -616 597
rect -682 547 -666 581
rect -632 547 -616 581
rect -682 531 -616 547
rect -564 581 -498 597
rect -564 547 -548 581
rect -514 547 -498 581
rect -564 531 -498 547
rect -446 581 -380 597
rect -446 547 -430 581
rect -396 547 -380 581
rect -446 531 -380 547
rect -328 581 -262 597
rect -328 547 -312 581
rect -278 547 -262 581
rect -328 531 -262 547
rect -210 581 -144 597
rect -210 547 -194 581
rect -160 547 -144 581
rect -210 531 -144 547
rect -92 581 -26 597
rect -92 547 -76 581
rect -42 547 -26 581
rect -92 531 -26 547
rect 26 581 92 597
rect 26 547 42 581
rect 76 547 92 581
rect 26 531 92 547
rect 144 581 210 597
rect 144 547 160 581
rect 194 547 210 581
rect 144 531 210 547
rect 262 581 328 597
rect 262 547 278 581
rect 312 547 328 581
rect 262 531 328 547
rect 380 581 446 597
rect 380 547 396 581
rect 430 547 446 581
rect 380 531 446 547
rect 498 581 564 597
rect 498 547 514 581
rect 548 547 564 581
rect 498 531 564 547
rect 616 581 682 597
rect 616 547 632 581
rect 666 547 682 581
rect 616 531 682 547
rect -679 509 -619 531
rect -561 509 -501 531
rect -443 509 -383 531
rect -325 509 -265 531
rect -207 509 -147 531
rect -89 509 -29 531
rect 29 509 89 531
rect 147 509 207 531
rect 265 509 325 531
rect 383 509 443 531
rect 501 509 561 531
rect 619 509 679 531
rect -679 87 -619 109
rect -561 87 -501 109
rect -443 87 -383 109
rect -325 87 -265 109
rect -207 87 -147 109
rect -89 87 -29 109
rect 29 87 89 109
rect 147 87 207 109
rect 265 87 325 109
rect 383 87 443 109
rect 501 87 561 109
rect 619 87 679 109
rect -682 71 -616 87
rect -682 37 -666 71
rect -632 37 -616 71
rect -682 21 -616 37
rect -564 71 -498 87
rect -564 37 -548 71
rect -514 37 -498 71
rect -564 21 -498 37
rect -446 71 -380 87
rect -446 37 -430 71
rect -396 37 -380 71
rect -446 21 -380 37
rect -328 71 -262 87
rect -328 37 -312 71
rect -278 37 -262 71
rect -328 21 -262 37
rect -210 71 -144 87
rect -210 37 -194 71
rect -160 37 -144 71
rect -210 21 -144 37
rect -92 71 -26 87
rect -92 37 -76 71
rect -42 37 -26 71
rect -92 21 -26 37
rect 26 71 92 87
rect 26 37 42 71
rect 76 37 92 71
rect 26 21 92 37
rect 144 71 210 87
rect 144 37 160 71
rect 194 37 210 71
rect 144 21 210 37
rect 262 71 328 87
rect 262 37 278 71
rect 312 37 328 71
rect 262 21 328 37
rect 380 71 446 87
rect 380 37 396 71
rect 430 37 446 71
rect 380 21 446 37
rect 498 71 564 87
rect 498 37 514 71
rect 548 37 564 71
rect 498 21 564 37
rect 616 71 682 87
rect 616 37 632 71
rect 666 37 682 71
rect 616 21 682 37
rect -682 -37 -616 -21
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -682 -87 -616 -71
rect -564 -37 -498 -21
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -564 -87 -498 -71
rect -446 -37 -380 -21
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -446 -87 -380 -71
rect -328 -37 -262 -21
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -328 -87 -262 -71
rect -210 -37 -144 -21
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -210 -87 -144 -71
rect -92 -37 -26 -21
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect -92 -87 -26 -71
rect 26 -37 92 -21
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 26 -87 92 -71
rect 144 -37 210 -21
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 144 -87 210 -71
rect 262 -37 328 -21
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 262 -87 328 -71
rect 380 -37 446 -21
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 380 -87 446 -71
rect 498 -37 564 -21
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 498 -87 564 -71
rect 616 -37 682 -21
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 616 -87 682 -71
rect -679 -109 -619 -87
rect -561 -109 -501 -87
rect -443 -109 -383 -87
rect -325 -109 -265 -87
rect -207 -109 -147 -87
rect -89 -109 -29 -87
rect 29 -109 89 -87
rect 147 -109 207 -87
rect 265 -109 325 -87
rect 383 -109 443 -87
rect 501 -109 561 -87
rect 619 -109 679 -87
rect -679 -531 -619 -509
rect -561 -531 -501 -509
rect -443 -531 -383 -509
rect -325 -531 -265 -509
rect -207 -531 -147 -509
rect -89 -531 -29 -509
rect 29 -531 89 -509
rect 147 -531 207 -509
rect 265 -531 325 -509
rect 383 -531 443 -509
rect 501 -531 561 -509
rect 619 -531 679 -509
rect -682 -547 -616 -531
rect -682 -581 -666 -547
rect -632 -581 -616 -547
rect -682 -597 -616 -581
rect -564 -547 -498 -531
rect -564 -581 -548 -547
rect -514 -581 -498 -547
rect -564 -597 -498 -581
rect -446 -547 -380 -531
rect -446 -581 -430 -547
rect -396 -581 -380 -547
rect -446 -597 -380 -581
rect -328 -547 -262 -531
rect -328 -581 -312 -547
rect -278 -581 -262 -547
rect -328 -597 -262 -581
rect -210 -547 -144 -531
rect -210 -581 -194 -547
rect -160 -581 -144 -547
rect -210 -597 -144 -581
rect -92 -547 -26 -531
rect -92 -581 -76 -547
rect -42 -581 -26 -547
rect -92 -597 -26 -581
rect 26 -547 92 -531
rect 26 -581 42 -547
rect 76 -581 92 -547
rect 26 -597 92 -581
rect 144 -547 210 -531
rect 144 -581 160 -547
rect 194 -581 210 -547
rect 144 -597 210 -581
rect 262 -547 328 -531
rect 262 -581 278 -547
rect 312 -581 328 -547
rect 262 -597 328 -581
rect 380 -547 446 -531
rect 380 -581 396 -547
rect 430 -581 446 -547
rect 380 -597 446 -581
rect 498 -547 564 -531
rect 498 -581 514 -547
rect 548 -581 564 -547
rect 498 -597 564 -581
rect 616 -547 682 -531
rect 616 -581 632 -547
rect 666 -581 682 -547
rect 616 -597 682 -581
<< polycont >>
rect -666 547 -632 581
rect -548 547 -514 581
rect -430 547 -396 581
rect -312 547 -278 581
rect -194 547 -160 581
rect -76 547 -42 581
rect 42 547 76 581
rect 160 547 194 581
rect 278 547 312 581
rect 396 547 430 581
rect 514 547 548 581
rect 632 547 666 581
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect -666 -581 -632 -547
rect -548 -581 -514 -547
rect -430 -581 -396 -547
rect -312 -581 -278 -547
rect -194 -581 -160 -547
rect -76 -581 -42 -547
rect 42 -581 76 -547
rect 160 -581 194 -547
rect 278 -581 312 -547
rect 396 -581 430 -547
rect 514 -581 548 -547
rect 632 -581 666 -547
<< locali >>
rect -839 649 -743 683
rect 743 649 839 683
rect -839 587 -805 649
rect 805 587 839 649
rect -682 547 -666 581
rect -632 547 -616 581
rect -564 547 -548 581
rect -514 547 -498 581
rect -446 547 -430 581
rect -396 547 -380 581
rect -328 547 -312 581
rect -278 547 -262 581
rect -210 547 -194 581
rect -160 547 -144 581
rect -92 547 -76 581
rect -42 547 -26 581
rect 26 547 42 581
rect 76 547 92 581
rect 144 547 160 581
rect 194 547 210 581
rect 262 547 278 581
rect 312 547 328 581
rect 380 547 396 581
rect 430 547 446 581
rect 498 547 514 581
rect 548 547 564 581
rect 616 547 632 581
rect 666 547 682 581
rect -725 497 -691 513
rect -725 105 -691 121
rect -607 497 -573 513
rect -607 105 -573 121
rect -489 497 -455 513
rect -489 105 -455 121
rect -371 497 -337 513
rect -371 105 -337 121
rect -253 497 -219 513
rect -253 105 -219 121
rect -135 497 -101 513
rect -135 105 -101 121
rect -17 497 17 513
rect -17 105 17 121
rect 101 497 135 513
rect 101 105 135 121
rect 219 497 253 513
rect 219 105 253 121
rect 337 497 371 513
rect 337 105 371 121
rect 455 497 489 513
rect 455 105 489 121
rect 573 497 607 513
rect 573 105 607 121
rect 691 497 725 513
rect 691 105 725 121
rect -682 37 -666 71
rect -632 37 -616 71
rect -564 37 -548 71
rect -514 37 -498 71
rect -446 37 -430 71
rect -396 37 -380 71
rect -328 37 -312 71
rect -278 37 -262 71
rect -210 37 -194 71
rect -160 37 -144 71
rect -92 37 -76 71
rect -42 37 -26 71
rect 26 37 42 71
rect 76 37 92 71
rect 144 37 160 71
rect 194 37 210 71
rect 262 37 278 71
rect 312 37 328 71
rect 380 37 396 71
rect 430 37 446 71
rect 498 37 514 71
rect 548 37 564 71
rect 616 37 632 71
rect 666 37 682 71
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 616 -71 632 -37
rect 666 -71 682 -37
rect -725 -121 -691 -105
rect -725 -513 -691 -497
rect -607 -121 -573 -105
rect -607 -513 -573 -497
rect -489 -121 -455 -105
rect -489 -513 -455 -497
rect -371 -121 -337 -105
rect -371 -513 -337 -497
rect -253 -121 -219 -105
rect -253 -513 -219 -497
rect -135 -121 -101 -105
rect -135 -513 -101 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 101 -121 135 -105
rect 101 -513 135 -497
rect 219 -121 253 -105
rect 219 -513 253 -497
rect 337 -121 371 -105
rect 337 -513 371 -497
rect 455 -121 489 -105
rect 455 -513 489 -497
rect 573 -121 607 -105
rect 573 -513 607 -497
rect 691 -121 725 -105
rect 691 -513 725 -497
rect -682 -581 -666 -547
rect -632 -581 -616 -547
rect -564 -581 -548 -547
rect -514 -581 -498 -547
rect -446 -581 -430 -547
rect -396 -581 -380 -547
rect -328 -581 -312 -547
rect -278 -581 -262 -547
rect -210 -581 -194 -547
rect -160 -581 -144 -547
rect -92 -581 -76 -547
rect -42 -581 -26 -547
rect 26 -581 42 -547
rect 76 -581 92 -547
rect 144 -581 160 -547
rect 194 -581 210 -547
rect 262 -581 278 -547
rect 312 -581 328 -547
rect 380 -581 396 -547
rect 430 -581 446 -547
rect 498 -581 514 -547
rect 548 -581 564 -547
rect 616 -581 632 -547
rect 666 -581 682 -547
rect -839 -649 -805 -587
rect 805 -649 839 -587
rect -839 -683 -743 -649
rect 743 -683 839 -649
<< viali >>
rect -666 547 -632 581
rect -548 547 -514 581
rect -430 547 -396 581
rect -312 547 -278 581
rect -194 547 -160 581
rect -76 547 -42 581
rect 42 547 76 581
rect 160 547 194 581
rect 278 547 312 581
rect 396 547 430 581
rect 514 547 548 581
rect 632 547 666 581
rect -725 121 -691 497
rect -607 121 -573 497
rect -489 121 -455 497
rect -371 121 -337 497
rect -253 121 -219 497
rect -135 121 -101 497
rect -17 121 17 497
rect 101 121 135 497
rect 219 121 253 497
rect 337 121 371 497
rect 455 121 489 497
rect 573 121 607 497
rect 691 121 725 497
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect -725 -497 -691 -121
rect -607 -497 -573 -121
rect -489 -497 -455 -121
rect -371 -497 -337 -121
rect -253 -497 -219 -121
rect -135 -497 -101 -121
rect -17 -497 17 -121
rect 101 -497 135 -121
rect 219 -497 253 -121
rect 337 -497 371 -121
rect 455 -497 489 -121
rect 573 -497 607 -121
rect 691 -497 725 -121
rect -666 -581 -632 -547
rect -548 -581 -514 -547
rect -430 -581 -396 -547
rect -312 -581 -278 -547
rect -194 -581 -160 -547
rect -76 -581 -42 -547
rect 42 -581 76 -547
rect 160 -581 194 -547
rect 278 -581 312 -547
rect 396 -581 430 -547
rect 514 -581 548 -547
rect 632 -581 666 -547
<< metal1 >>
rect -678 581 -620 587
rect -678 547 -666 581
rect -632 547 -620 581
rect -678 541 -620 547
rect -560 581 -502 587
rect -560 547 -548 581
rect -514 547 -502 581
rect -560 541 -502 547
rect -442 581 -384 587
rect -442 547 -430 581
rect -396 547 -384 581
rect -442 541 -384 547
rect -324 581 -266 587
rect -324 547 -312 581
rect -278 547 -266 581
rect -324 541 -266 547
rect -206 581 -148 587
rect -206 547 -194 581
rect -160 547 -148 581
rect -206 541 -148 547
rect -88 581 -30 587
rect -88 547 -76 581
rect -42 547 -30 581
rect -88 541 -30 547
rect 30 581 88 587
rect 30 547 42 581
rect 76 547 88 581
rect 30 541 88 547
rect 148 581 206 587
rect 148 547 160 581
rect 194 547 206 581
rect 148 541 206 547
rect 266 581 324 587
rect 266 547 278 581
rect 312 547 324 581
rect 266 541 324 547
rect 384 581 442 587
rect 384 547 396 581
rect 430 547 442 581
rect 384 541 442 547
rect 502 581 560 587
rect 502 547 514 581
rect 548 547 560 581
rect 502 541 560 547
rect 620 581 678 587
rect 620 547 632 581
rect 666 547 678 581
rect 620 541 678 547
rect -731 497 -685 509
rect -731 121 -725 497
rect -691 121 -685 497
rect -731 109 -685 121
rect -613 497 -567 509
rect -613 121 -607 497
rect -573 121 -567 497
rect -613 109 -567 121
rect -495 497 -449 509
rect -495 121 -489 497
rect -455 121 -449 497
rect -495 109 -449 121
rect -377 497 -331 509
rect -377 121 -371 497
rect -337 121 -331 497
rect -377 109 -331 121
rect -259 497 -213 509
rect -259 121 -253 497
rect -219 121 -213 497
rect -259 109 -213 121
rect -141 497 -95 509
rect -141 121 -135 497
rect -101 121 -95 497
rect -141 109 -95 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 95 497 141 509
rect 95 121 101 497
rect 135 121 141 497
rect 95 109 141 121
rect 213 497 259 509
rect 213 121 219 497
rect 253 121 259 497
rect 213 109 259 121
rect 331 497 377 509
rect 331 121 337 497
rect 371 121 377 497
rect 331 109 377 121
rect 449 497 495 509
rect 449 121 455 497
rect 489 121 495 497
rect 449 109 495 121
rect 567 497 613 509
rect 567 121 573 497
rect 607 121 613 497
rect 567 109 613 121
rect 685 497 731 509
rect 685 121 691 497
rect 725 121 731 497
rect 685 109 731 121
rect -678 71 -620 77
rect -678 37 -666 71
rect -632 37 -620 71
rect -678 31 -620 37
rect -560 71 -502 77
rect -560 37 -548 71
rect -514 37 -502 71
rect -560 31 -502 37
rect -442 71 -384 77
rect -442 37 -430 71
rect -396 37 -384 71
rect -442 31 -384 37
rect -324 71 -266 77
rect -324 37 -312 71
rect -278 37 -266 71
rect -324 31 -266 37
rect -206 71 -148 77
rect -206 37 -194 71
rect -160 37 -148 71
rect -206 31 -148 37
rect -88 71 -30 77
rect -88 37 -76 71
rect -42 37 -30 71
rect -88 31 -30 37
rect 30 71 88 77
rect 30 37 42 71
rect 76 37 88 71
rect 30 31 88 37
rect 148 71 206 77
rect 148 37 160 71
rect 194 37 206 71
rect 148 31 206 37
rect 266 71 324 77
rect 266 37 278 71
rect 312 37 324 71
rect 266 31 324 37
rect 384 71 442 77
rect 384 37 396 71
rect 430 37 442 71
rect 384 31 442 37
rect 502 71 560 77
rect 502 37 514 71
rect 548 37 560 71
rect 502 31 560 37
rect 620 71 678 77
rect 620 37 632 71
rect 666 37 678 71
rect 620 31 678 37
rect -678 -37 -620 -31
rect -678 -71 -666 -37
rect -632 -71 -620 -37
rect -678 -77 -620 -71
rect -560 -37 -502 -31
rect -560 -71 -548 -37
rect -514 -71 -502 -37
rect -560 -77 -502 -71
rect -442 -37 -384 -31
rect -442 -71 -430 -37
rect -396 -71 -384 -37
rect -442 -77 -384 -71
rect -324 -37 -266 -31
rect -324 -71 -312 -37
rect -278 -71 -266 -37
rect -324 -77 -266 -71
rect -206 -37 -148 -31
rect -206 -71 -194 -37
rect -160 -71 -148 -37
rect -206 -77 -148 -71
rect -88 -37 -30 -31
rect -88 -71 -76 -37
rect -42 -71 -30 -37
rect -88 -77 -30 -71
rect 30 -37 88 -31
rect 30 -71 42 -37
rect 76 -71 88 -37
rect 30 -77 88 -71
rect 148 -37 206 -31
rect 148 -71 160 -37
rect 194 -71 206 -37
rect 148 -77 206 -71
rect 266 -37 324 -31
rect 266 -71 278 -37
rect 312 -71 324 -37
rect 266 -77 324 -71
rect 384 -37 442 -31
rect 384 -71 396 -37
rect 430 -71 442 -37
rect 384 -77 442 -71
rect 502 -37 560 -31
rect 502 -71 514 -37
rect 548 -71 560 -37
rect 502 -77 560 -71
rect 620 -37 678 -31
rect 620 -71 632 -37
rect 666 -71 678 -37
rect 620 -77 678 -71
rect -731 -121 -685 -109
rect -731 -497 -725 -121
rect -691 -497 -685 -121
rect -731 -509 -685 -497
rect -613 -121 -567 -109
rect -613 -497 -607 -121
rect -573 -497 -567 -121
rect -613 -509 -567 -497
rect -495 -121 -449 -109
rect -495 -497 -489 -121
rect -455 -497 -449 -121
rect -495 -509 -449 -497
rect -377 -121 -331 -109
rect -377 -497 -371 -121
rect -337 -497 -331 -121
rect -377 -509 -331 -497
rect -259 -121 -213 -109
rect -259 -497 -253 -121
rect -219 -497 -213 -121
rect -259 -509 -213 -497
rect -141 -121 -95 -109
rect -141 -497 -135 -121
rect -101 -497 -95 -121
rect -141 -509 -95 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 95 -121 141 -109
rect 95 -497 101 -121
rect 135 -497 141 -121
rect 95 -509 141 -497
rect 213 -121 259 -109
rect 213 -497 219 -121
rect 253 -497 259 -121
rect 213 -509 259 -497
rect 331 -121 377 -109
rect 331 -497 337 -121
rect 371 -497 377 -121
rect 331 -509 377 -497
rect 449 -121 495 -109
rect 449 -497 455 -121
rect 489 -497 495 -121
rect 449 -509 495 -497
rect 567 -121 613 -109
rect 567 -497 573 -121
rect 607 -497 613 -121
rect 567 -509 613 -497
rect 685 -121 731 -109
rect 685 -497 691 -121
rect 725 -497 731 -121
rect 685 -509 731 -497
rect -678 -547 -620 -541
rect -678 -581 -666 -547
rect -632 -581 -620 -547
rect -678 -587 -620 -581
rect -560 -547 -502 -541
rect -560 -581 -548 -547
rect -514 -581 -502 -547
rect -560 -587 -502 -581
rect -442 -547 -384 -541
rect -442 -581 -430 -547
rect -396 -581 -384 -547
rect -442 -587 -384 -581
rect -324 -547 -266 -541
rect -324 -581 -312 -547
rect -278 -581 -266 -547
rect -324 -587 -266 -581
rect -206 -547 -148 -541
rect -206 -581 -194 -547
rect -160 -581 -148 -547
rect -206 -587 -148 -581
rect -88 -547 -30 -541
rect -88 -581 -76 -547
rect -42 -581 -30 -547
rect -88 -587 -30 -581
rect 30 -547 88 -541
rect 30 -581 42 -547
rect 76 -581 88 -547
rect 30 -587 88 -581
rect 148 -547 206 -541
rect 148 -581 160 -547
rect 194 -581 206 -547
rect 148 -587 206 -581
rect 266 -547 324 -541
rect 266 -581 278 -547
rect 312 -581 324 -547
rect 266 -587 324 -581
rect 384 -547 442 -541
rect 384 -581 396 -547
rect 430 -581 442 -547
rect 384 -587 442 -581
rect 502 -547 560 -541
rect 502 -581 514 -547
rect 548 -581 560 -547
rect 502 -587 560 -581
rect 620 -547 678 -541
rect 620 -581 632 -547
rect 666 -581 678 -547
rect 620 -587 678 -581
<< properties >>
string FIXED_BBOX -822 -666 822 666
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.3 m 2 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
