magic
tech sky130B
magscale 1 2
timestamp 1653911185
<< metal4 >>
rect -2351 3059 2351 3100
rect -2351 -3059 2095 3059
rect 2331 -3059 2351 3059
rect -2351 -3100 2351 -3059
<< via4 >>
rect 2095 -3059 2331 3059
<< mimcap2 >>
rect -2251 2960 1749 3000
rect -2251 -2960 -2211 2960
rect 1709 -2960 1749 2960
rect -2251 -3000 1749 -2960
<< mimcap2contact >>
rect -2211 -2960 1709 2960
<< metal5 >>
rect 2053 3059 2373 3101
rect -2235 2960 1733 2984
rect -2235 -2960 -2211 2960
rect 1709 -2960 1733 2960
rect -2235 -2984 1733 -2960
rect 2053 -3059 2095 3059
rect 2331 -3059 2373 3059
rect 2053 -3101 2373 -3059
<< properties >>
string FIXED_BBOX -2351 -3100 1849 3100
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20 l 30 val 1.219k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
