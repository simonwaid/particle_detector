magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< error_p >>
rect -557 1199 -499 1205
rect -365 1199 -307 1205
rect -173 1199 -115 1205
rect 19 1199 77 1205
rect 211 1199 269 1205
rect 403 1199 461 1205
rect -557 1165 -545 1199
rect -365 1165 -353 1199
rect -173 1165 -161 1199
rect 19 1165 31 1199
rect 211 1165 223 1199
rect 403 1165 415 1199
rect -557 1159 -499 1165
rect -365 1159 -307 1165
rect -173 1159 -115 1165
rect 19 1159 77 1165
rect 211 1159 269 1165
rect 403 1159 461 1165
rect -461 689 -403 695
rect -269 689 -211 695
rect -77 689 -19 695
rect 115 689 173 695
rect 307 689 365 695
rect 499 689 557 695
rect -461 655 -449 689
rect -269 655 -257 689
rect -77 655 -65 689
rect 115 655 127 689
rect 307 655 319 689
rect 499 655 511 689
rect -461 649 -403 655
rect -269 649 -211 655
rect -77 649 -19 655
rect 115 649 173 655
rect 307 649 365 655
rect 499 649 557 655
rect -461 581 -403 587
rect -269 581 -211 587
rect -77 581 -19 587
rect 115 581 173 587
rect 307 581 365 587
rect 499 581 557 587
rect -461 547 -449 581
rect -269 547 -257 581
rect -77 547 -65 581
rect 115 547 127 581
rect 307 547 319 581
rect 499 547 511 581
rect -461 541 -403 547
rect -269 541 -211 547
rect -77 541 -19 547
rect 115 541 173 547
rect 307 541 365 547
rect 499 541 557 547
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect -461 -547 -403 -541
rect -269 -547 -211 -541
rect -77 -547 -19 -541
rect 115 -547 173 -541
rect 307 -547 365 -541
rect 499 -547 557 -541
rect -461 -581 -449 -547
rect -269 -581 -257 -547
rect -77 -581 -65 -547
rect 115 -581 127 -547
rect 307 -581 319 -547
rect 499 -581 511 -547
rect -461 -587 -403 -581
rect -269 -587 -211 -581
rect -77 -587 -19 -581
rect 115 -587 173 -581
rect 307 -587 365 -581
rect 499 -587 557 -581
rect -461 -655 -403 -649
rect -269 -655 -211 -649
rect -77 -655 -19 -649
rect 115 -655 173 -649
rect 307 -655 365 -649
rect 499 -655 557 -649
rect -461 -689 -449 -655
rect -269 -689 -257 -655
rect -77 -689 -65 -655
rect 115 -689 127 -655
rect 307 -689 319 -655
rect 499 -689 511 -655
rect -461 -695 -403 -689
rect -269 -695 -211 -689
rect -77 -695 -19 -689
rect 115 -695 173 -689
rect 307 -695 365 -689
rect 499 -695 557 -689
rect -557 -1165 -499 -1159
rect -365 -1165 -307 -1159
rect -173 -1165 -115 -1159
rect 19 -1165 77 -1159
rect 211 -1165 269 -1159
rect 403 -1165 461 -1159
rect -557 -1199 -545 -1165
rect -365 -1199 -353 -1165
rect -173 -1199 -161 -1165
rect 19 -1199 31 -1165
rect 211 -1199 223 -1165
rect 403 -1199 415 -1165
rect -557 -1205 -499 -1199
rect -365 -1205 -307 -1199
rect -173 -1205 -115 -1199
rect 19 -1205 77 -1199
rect 211 -1205 269 -1199
rect 403 -1205 461 -1199
<< pwell >>
rect -743 -1337 743 1337
<< nmos >>
rect -543 727 -513 1127
rect -447 727 -417 1127
rect -351 727 -321 1127
rect -255 727 -225 1127
rect -159 727 -129 1127
rect -63 727 -33 1127
rect 33 727 63 1127
rect 129 727 159 1127
rect 225 727 255 1127
rect 321 727 351 1127
rect 417 727 447 1127
rect 513 727 543 1127
rect -543 109 -513 509
rect -447 109 -417 509
rect -351 109 -321 509
rect -255 109 -225 509
rect -159 109 -129 509
rect -63 109 -33 509
rect 33 109 63 509
rect 129 109 159 509
rect 225 109 255 509
rect 321 109 351 509
rect 417 109 447 509
rect 513 109 543 509
rect -543 -509 -513 -109
rect -447 -509 -417 -109
rect -351 -509 -321 -109
rect -255 -509 -225 -109
rect -159 -509 -129 -109
rect -63 -509 -33 -109
rect 33 -509 63 -109
rect 129 -509 159 -109
rect 225 -509 255 -109
rect 321 -509 351 -109
rect 417 -509 447 -109
rect 513 -509 543 -109
rect -543 -1127 -513 -727
rect -447 -1127 -417 -727
rect -351 -1127 -321 -727
rect -255 -1127 -225 -727
rect -159 -1127 -129 -727
rect -63 -1127 -33 -727
rect 33 -1127 63 -727
rect 129 -1127 159 -727
rect 225 -1127 255 -727
rect 321 -1127 351 -727
rect 417 -1127 447 -727
rect 513 -1127 543 -727
<< ndiff >>
rect -605 1115 -543 1127
rect -605 739 -593 1115
rect -559 739 -543 1115
rect -605 727 -543 739
rect -513 1115 -447 1127
rect -513 739 -497 1115
rect -463 739 -447 1115
rect -513 727 -447 739
rect -417 1115 -351 1127
rect -417 739 -401 1115
rect -367 739 -351 1115
rect -417 727 -351 739
rect -321 1115 -255 1127
rect -321 739 -305 1115
rect -271 739 -255 1115
rect -321 727 -255 739
rect -225 1115 -159 1127
rect -225 739 -209 1115
rect -175 739 -159 1115
rect -225 727 -159 739
rect -129 1115 -63 1127
rect -129 739 -113 1115
rect -79 739 -63 1115
rect -129 727 -63 739
rect -33 1115 33 1127
rect -33 739 -17 1115
rect 17 739 33 1115
rect -33 727 33 739
rect 63 1115 129 1127
rect 63 739 79 1115
rect 113 739 129 1115
rect 63 727 129 739
rect 159 1115 225 1127
rect 159 739 175 1115
rect 209 739 225 1115
rect 159 727 225 739
rect 255 1115 321 1127
rect 255 739 271 1115
rect 305 739 321 1115
rect 255 727 321 739
rect 351 1115 417 1127
rect 351 739 367 1115
rect 401 739 417 1115
rect 351 727 417 739
rect 447 1115 513 1127
rect 447 739 463 1115
rect 497 739 513 1115
rect 447 727 513 739
rect 543 1115 605 1127
rect 543 739 559 1115
rect 593 739 605 1115
rect 543 727 605 739
rect -605 497 -543 509
rect -605 121 -593 497
rect -559 121 -543 497
rect -605 109 -543 121
rect -513 497 -447 509
rect -513 121 -497 497
rect -463 121 -447 497
rect -513 109 -447 121
rect -417 497 -351 509
rect -417 121 -401 497
rect -367 121 -351 497
rect -417 109 -351 121
rect -321 497 -255 509
rect -321 121 -305 497
rect -271 121 -255 497
rect -321 109 -255 121
rect -225 497 -159 509
rect -225 121 -209 497
rect -175 121 -159 497
rect -225 109 -159 121
rect -129 497 -63 509
rect -129 121 -113 497
rect -79 121 -63 497
rect -129 109 -63 121
rect -33 497 33 509
rect -33 121 -17 497
rect 17 121 33 497
rect -33 109 33 121
rect 63 497 129 509
rect 63 121 79 497
rect 113 121 129 497
rect 63 109 129 121
rect 159 497 225 509
rect 159 121 175 497
rect 209 121 225 497
rect 159 109 225 121
rect 255 497 321 509
rect 255 121 271 497
rect 305 121 321 497
rect 255 109 321 121
rect 351 497 417 509
rect 351 121 367 497
rect 401 121 417 497
rect 351 109 417 121
rect 447 497 513 509
rect 447 121 463 497
rect 497 121 513 497
rect 447 109 513 121
rect 543 497 605 509
rect 543 121 559 497
rect 593 121 605 497
rect 543 109 605 121
rect -605 -121 -543 -109
rect -605 -497 -593 -121
rect -559 -497 -543 -121
rect -605 -509 -543 -497
rect -513 -121 -447 -109
rect -513 -497 -497 -121
rect -463 -497 -447 -121
rect -513 -509 -447 -497
rect -417 -121 -351 -109
rect -417 -497 -401 -121
rect -367 -497 -351 -121
rect -417 -509 -351 -497
rect -321 -121 -255 -109
rect -321 -497 -305 -121
rect -271 -497 -255 -121
rect -321 -509 -255 -497
rect -225 -121 -159 -109
rect -225 -497 -209 -121
rect -175 -497 -159 -121
rect -225 -509 -159 -497
rect -129 -121 -63 -109
rect -129 -497 -113 -121
rect -79 -497 -63 -121
rect -129 -509 -63 -497
rect -33 -121 33 -109
rect -33 -497 -17 -121
rect 17 -497 33 -121
rect -33 -509 33 -497
rect 63 -121 129 -109
rect 63 -497 79 -121
rect 113 -497 129 -121
rect 63 -509 129 -497
rect 159 -121 225 -109
rect 159 -497 175 -121
rect 209 -497 225 -121
rect 159 -509 225 -497
rect 255 -121 321 -109
rect 255 -497 271 -121
rect 305 -497 321 -121
rect 255 -509 321 -497
rect 351 -121 417 -109
rect 351 -497 367 -121
rect 401 -497 417 -121
rect 351 -509 417 -497
rect 447 -121 513 -109
rect 447 -497 463 -121
rect 497 -497 513 -121
rect 447 -509 513 -497
rect 543 -121 605 -109
rect 543 -497 559 -121
rect 593 -497 605 -121
rect 543 -509 605 -497
rect -605 -739 -543 -727
rect -605 -1115 -593 -739
rect -559 -1115 -543 -739
rect -605 -1127 -543 -1115
rect -513 -739 -447 -727
rect -513 -1115 -497 -739
rect -463 -1115 -447 -739
rect -513 -1127 -447 -1115
rect -417 -739 -351 -727
rect -417 -1115 -401 -739
rect -367 -1115 -351 -739
rect -417 -1127 -351 -1115
rect -321 -739 -255 -727
rect -321 -1115 -305 -739
rect -271 -1115 -255 -739
rect -321 -1127 -255 -1115
rect -225 -739 -159 -727
rect -225 -1115 -209 -739
rect -175 -1115 -159 -739
rect -225 -1127 -159 -1115
rect -129 -739 -63 -727
rect -129 -1115 -113 -739
rect -79 -1115 -63 -739
rect -129 -1127 -63 -1115
rect -33 -739 33 -727
rect -33 -1115 -17 -739
rect 17 -1115 33 -739
rect -33 -1127 33 -1115
rect 63 -739 129 -727
rect 63 -1115 79 -739
rect 113 -1115 129 -739
rect 63 -1127 129 -1115
rect 159 -739 225 -727
rect 159 -1115 175 -739
rect 209 -1115 225 -739
rect 159 -1127 225 -1115
rect 255 -739 321 -727
rect 255 -1115 271 -739
rect 305 -1115 321 -739
rect 255 -1127 321 -1115
rect 351 -739 417 -727
rect 351 -1115 367 -739
rect 401 -1115 417 -739
rect 351 -1127 417 -1115
rect 447 -739 513 -727
rect 447 -1115 463 -739
rect 497 -1115 513 -739
rect 447 -1127 513 -1115
rect 543 -739 605 -727
rect 543 -1115 559 -739
rect 593 -1115 605 -739
rect 543 -1127 605 -1115
<< ndiffc >>
rect -593 739 -559 1115
rect -497 739 -463 1115
rect -401 739 -367 1115
rect -305 739 -271 1115
rect -209 739 -175 1115
rect -113 739 -79 1115
rect -17 739 17 1115
rect 79 739 113 1115
rect 175 739 209 1115
rect 271 739 305 1115
rect 367 739 401 1115
rect 463 739 497 1115
rect 559 739 593 1115
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect -593 -1115 -559 -739
rect -497 -1115 -463 -739
rect -401 -1115 -367 -739
rect -305 -1115 -271 -739
rect -209 -1115 -175 -739
rect -113 -1115 -79 -739
rect -17 -1115 17 -739
rect 79 -1115 113 -739
rect 175 -1115 209 -739
rect 271 -1115 305 -739
rect 367 -1115 401 -739
rect 463 -1115 497 -739
rect 559 -1115 593 -739
<< psubdiff >>
rect -707 1267 -611 1301
rect 611 1267 707 1301
rect -707 1205 -673 1267
rect 673 1205 707 1267
rect -707 -1267 -673 -1205
rect 673 -1267 707 -1205
rect -707 -1301 -611 -1267
rect 611 -1301 707 -1267
<< psubdiffcont >>
rect -611 1267 611 1301
rect -707 -1205 -673 1205
rect 673 -1205 707 1205
rect -611 -1301 611 -1267
<< poly >>
rect -561 1199 -495 1215
rect -561 1165 -545 1199
rect -511 1165 -495 1199
rect -561 1149 -495 1165
rect -369 1199 -303 1215
rect -369 1165 -353 1199
rect -319 1165 -303 1199
rect -543 1127 -513 1149
rect -447 1127 -417 1153
rect -369 1149 -303 1165
rect -177 1199 -111 1215
rect -177 1165 -161 1199
rect -127 1165 -111 1199
rect -351 1127 -321 1149
rect -255 1127 -225 1153
rect -177 1149 -111 1165
rect 15 1199 81 1215
rect 15 1165 31 1199
rect 65 1165 81 1199
rect -159 1127 -129 1149
rect -63 1127 -33 1153
rect 15 1149 81 1165
rect 207 1199 273 1215
rect 207 1165 223 1199
rect 257 1165 273 1199
rect 33 1127 63 1149
rect 129 1127 159 1153
rect 207 1149 273 1165
rect 399 1199 465 1215
rect 399 1165 415 1199
rect 449 1165 465 1199
rect 225 1127 255 1149
rect 321 1127 351 1153
rect 399 1149 465 1165
rect 417 1127 447 1149
rect 513 1127 543 1153
rect -543 701 -513 727
rect -447 705 -417 727
rect -465 689 -399 705
rect -351 701 -321 727
rect -255 705 -225 727
rect -465 655 -449 689
rect -415 655 -399 689
rect -465 639 -399 655
rect -273 689 -207 705
rect -159 701 -129 727
rect -63 705 -33 727
rect -273 655 -257 689
rect -223 655 -207 689
rect -273 639 -207 655
rect -81 689 -15 705
rect 33 701 63 727
rect 129 705 159 727
rect -81 655 -65 689
rect -31 655 -15 689
rect -81 639 -15 655
rect 111 689 177 705
rect 225 701 255 727
rect 321 705 351 727
rect 111 655 127 689
rect 161 655 177 689
rect 111 639 177 655
rect 303 689 369 705
rect 417 701 447 727
rect 513 705 543 727
rect 303 655 319 689
rect 353 655 369 689
rect 303 639 369 655
rect 495 689 561 705
rect 495 655 511 689
rect 545 655 561 689
rect 495 639 561 655
rect -465 581 -399 597
rect -465 547 -449 581
rect -415 547 -399 581
rect -543 509 -513 535
rect -465 531 -399 547
rect -273 581 -207 597
rect -273 547 -257 581
rect -223 547 -207 581
rect -447 509 -417 531
rect -351 509 -321 535
rect -273 531 -207 547
rect -81 581 -15 597
rect -81 547 -65 581
rect -31 547 -15 581
rect -255 509 -225 531
rect -159 509 -129 535
rect -81 531 -15 547
rect 111 581 177 597
rect 111 547 127 581
rect 161 547 177 581
rect -63 509 -33 531
rect 33 509 63 535
rect 111 531 177 547
rect 303 581 369 597
rect 303 547 319 581
rect 353 547 369 581
rect 129 509 159 531
rect 225 509 255 535
rect 303 531 369 547
rect 495 581 561 597
rect 495 547 511 581
rect 545 547 561 581
rect 321 509 351 531
rect 417 509 447 535
rect 495 531 561 547
rect 513 509 543 531
rect -543 87 -513 109
rect -561 71 -495 87
rect -447 83 -417 109
rect -351 87 -321 109
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 513 83 543 109
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -543 -109 -513 -87
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 417 -109 447 -87
rect 513 -109 543 -83
rect -543 -535 -513 -509
rect -447 -531 -417 -509
rect -465 -547 -399 -531
rect -351 -535 -321 -509
rect -255 -531 -225 -509
rect -465 -581 -449 -547
rect -415 -581 -399 -547
rect -465 -597 -399 -581
rect -273 -547 -207 -531
rect -159 -535 -129 -509
rect -63 -531 -33 -509
rect -273 -581 -257 -547
rect -223 -581 -207 -547
rect -273 -597 -207 -581
rect -81 -547 -15 -531
rect 33 -535 63 -509
rect 129 -531 159 -509
rect -81 -581 -65 -547
rect -31 -581 -15 -547
rect -81 -597 -15 -581
rect 111 -547 177 -531
rect 225 -535 255 -509
rect 321 -531 351 -509
rect 111 -581 127 -547
rect 161 -581 177 -547
rect 111 -597 177 -581
rect 303 -547 369 -531
rect 417 -535 447 -509
rect 513 -531 543 -509
rect 303 -581 319 -547
rect 353 -581 369 -547
rect 303 -597 369 -581
rect 495 -547 561 -531
rect 495 -581 511 -547
rect 545 -581 561 -547
rect 495 -597 561 -581
rect -465 -655 -399 -639
rect -465 -689 -449 -655
rect -415 -689 -399 -655
rect -543 -727 -513 -701
rect -465 -705 -399 -689
rect -273 -655 -207 -639
rect -273 -689 -257 -655
rect -223 -689 -207 -655
rect -447 -727 -417 -705
rect -351 -727 -321 -701
rect -273 -705 -207 -689
rect -81 -655 -15 -639
rect -81 -689 -65 -655
rect -31 -689 -15 -655
rect -255 -727 -225 -705
rect -159 -727 -129 -701
rect -81 -705 -15 -689
rect 111 -655 177 -639
rect 111 -689 127 -655
rect 161 -689 177 -655
rect -63 -727 -33 -705
rect 33 -727 63 -701
rect 111 -705 177 -689
rect 303 -655 369 -639
rect 303 -689 319 -655
rect 353 -689 369 -655
rect 129 -727 159 -705
rect 225 -727 255 -701
rect 303 -705 369 -689
rect 495 -655 561 -639
rect 495 -689 511 -655
rect 545 -689 561 -655
rect 321 -727 351 -705
rect 417 -727 447 -701
rect 495 -705 561 -689
rect 513 -727 543 -705
rect -543 -1149 -513 -1127
rect -561 -1165 -495 -1149
rect -447 -1153 -417 -1127
rect -351 -1149 -321 -1127
rect -561 -1199 -545 -1165
rect -511 -1199 -495 -1165
rect -561 -1215 -495 -1199
rect -369 -1165 -303 -1149
rect -255 -1153 -225 -1127
rect -159 -1149 -129 -1127
rect -369 -1199 -353 -1165
rect -319 -1199 -303 -1165
rect -369 -1215 -303 -1199
rect -177 -1165 -111 -1149
rect -63 -1153 -33 -1127
rect 33 -1149 63 -1127
rect -177 -1199 -161 -1165
rect -127 -1199 -111 -1165
rect -177 -1215 -111 -1199
rect 15 -1165 81 -1149
rect 129 -1153 159 -1127
rect 225 -1149 255 -1127
rect 15 -1199 31 -1165
rect 65 -1199 81 -1165
rect 15 -1215 81 -1199
rect 207 -1165 273 -1149
rect 321 -1153 351 -1127
rect 417 -1149 447 -1127
rect 207 -1199 223 -1165
rect 257 -1199 273 -1165
rect 207 -1215 273 -1199
rect 399 -1165 465 -1149
rect 513 -1153 543 -1127
rect 399 -1199 415 -1165
rect 449 -1199 465 -1165
rect 399 -1215 465 -1199
<< polycont >>
rect -545 1165 -511 1199
rect -353 1165 -319 1199
rect -161 1165 -127 1199
rect 31 1165 65 1199
rect 223 1165 257 1199
rect 415 1165 449 1199
rect -449 655 -415 689
rect -257 655 -223 689
rect -65 655 -31 689
rect 127 655 161 689
rect 319 655 353 689
rect 511 655 545 689
rect -449 547 -415 581
rect -257 547 -223 581
rect -65 547 -31 581
rect 127 547 161 581
rect 319 547 353 581
rect 511 547 545 581
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -449 -581 -415 -547
rect -257 -581 -223 -547
rect -65 -581 -31 -547
rect 127 -581 161 -547
rect 319 -581 353 -547
rect 511 -581 545 -547
rect -449 -689 -415 -655
rect -257 -689 -223 -655
rect -65 -689 -31 -655
rect 127 -689 161 -655
rect 319 -689 353 -655
rect 511 -689 545 -655
rect -545 -1199 -511 -1165
rect -353 -1199 -319 -1165
rect -161 -1199 -127 -1165
rect 31 -1199 65 -1165
rect 223 -1199 257 -1165
rect 415 -1199 449 -1165
<< locali >>
rect -707 1267 -611 1301
rect 611 1267 707 1301
rect -707 1205 -673 1267
rect 673 1205 707 1267
rect -561 1165 -545 1199
rect -511 1165 -495 1199
rect -369 1165 -353 1199
rect -319 1165 -303 1199
rect -177 1165 -161 1199
rect -127 1165 -111 1199
rect 15 1165 31 1199
rect 65 1165 81 1199
rect 207 1165 223 1199
rect 257 1165 273 1199
rect 399 1165 415 1199
rect 449 1165 465 1199
rect -593 1115 -559 1131
rect -593 723 -559 739
rect -497 1115 -463 1131
rect -497 723 -463 739
rect -401 1115 -367 1131
rect -401 723 -367 739
rect -305 1115 -271 1131
rect -305 723 -271 739
rect -209 1115 -175 1131
rect -209 723 -175 739
rect -113 1115 -79 1131
rect -113 723 -79 739
rect -17 1115 17 1131
rect -17 723 17 739
rect 79 1115 113 1131
rect 79 723 113 739
rect 175 1115 209 1131
rect 175 723 209 739
rect 271 1115 305 1131
rect 271 723 305 739
rect 367 1115 401 1131
rect 367 723 401 739
rect 463 1115 497 1131
rect 463 723 497 739
rect 559 1115 593 1131
rect 559 723 593 739
rect -465 655 -449 689
rect -415 655 -399 689
rect -273 655 -257 689
rect -223 655 -207 689
rect -81 655 -65 689
rect -31 655 -15 689
rect 111 655 127 689
rect 161 655 177 689
rect 303 655 319 689
rect 353 655 369 689
rect 495 655 511 689
rect 545 655 561 689
rect -465 547 -449 581
rect -415 547 -399 581
rect -273 547 -257 581
rect -223 547 -207 581
rect -81 547 -65 581
rect -31 547 -15 581
rect 111 547 127 581
rect 161 547 177 581
rect 303 547 319 581
rect 353 547 369 581
rect 495 547 511 581
rect 545 547 561 581
rect -593 497 -559 513
rect -593 105 -559 121
rect -497 497 -463 513
rect -497 105 -463 121
rect -401 497 -367 513
rect -401 105 -367 121
rect -305 497 -271 513
rect -305 105 -271 121
rect -209 497 -175 513
rect -209 105 -175 121
rect -113 497 -79 513
rect -113 105 -79 121
rect -17 497 17 513
rect -17 105 17 121
rect 79 497 113 513
rect 79 105 113 121
rect 175 497 209 513
rect 175 105 209 121
rect 271 497 305 513
rect 271 105 305 121
rect 367 497 401 513
rect 367 105 401 121
rect 463 497 497 513
rect 463 105 497 121
rect 559 497 593 513
rect 559 105 593 121
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect -593 -121 -559 -105
rect -593 -513 -559 -497
rect -497 -121 -463 -105
rect -497 -513 -463 -497
rect -401 -121 -367 -105
rect -401 -513 -367 -497
rect -305 -121 -271 -105
rect -305 -513 -271 -497
rect -209 -121 -175 -105
rect -209 -513 -175 -497
rect -113 -121 -79 -105
rect -113 -513 -79 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 79 -121 113 -105
rect 79 -513 113 -497
rect 175 -121 209 -105
rect 175 -513 209 -497
rect 271 -121 305 -105
rect 271 -513 305 -497
rect 367 -121 401 -105
rect 367 -513 401 -497
rect 463 -121 497 -105
rect 463 -513 497 -497
rect 559 -121 593 -105
rect 559 -513 593 -497
rect -465 -581 -449 -547
rect -415 -581 -399 -547
rect -273 -581 -257 -547
rect -223 -581 -207 -547
rect -81 -581 -65 -547
rect -31 -581 -15 -547
rect 111 -581 127 -547
rect 161 -581 177 -547
rect 303 -581 319 -547
rect 353 -581 369 -547
rect 495 -581 511 -547
rect 545 -581 561 -547
rect -465 -689 -449 -655
rect -415 -689 -399 -655
rect -273 -689 -257 -655
rect -223 -689 -207 -655
rect -81 -689 -65 -655
rect -31 -689 -15 -655
rect 111 -689 127 -655
rect 161 -689 177 -655
rect 303 -689 319 -655
rect 353 -689 369 -655
rect 495 -689 511 -655
rect 545 -689 561 -655
rect -593 -739 -559 -723
rect -593 -1131 -559 -1115
rect -497 -739 -463 -723
rect -497 -1131 -463 -1115
rect -401 -739 -367 -723
rect -401 -1131 -367 -1115
rect -305 -739 -271 -723
rect -305 -1131 -271 -1115
rect -209 -739 -175 -723
rect -209 -1131 -175 -1115
rect -113 -739 -79 -723
rect -113 -1131 -79 -1115
rect -17 -739 17 -723
rect -17 -1131 17 -1115
rect 79 -739 113 -723
rect 79 -1131 113 -1115
rect 175 -739 209 -723
rect 175 -1131 209 -1115
rect 271 -739 305 -723
rect 271 -1131 305 -1115
rect 367 -739 401 -723
rect 367 -1131 401 -1115
rect 463 -739 497 -723
rect 463 -1131 497 -1115
rect 559 -739 593 -723
rect 559 -1131 593 -1115
rect -561 -1199 -545 -1165
rect -511 -1199 -495 -1165
rect -369 -1199 -353 -1165
rect -319 -1199 -303 -1165
rect -177 -1199 -161 -1165
rect -127 -1199 -111 -1165
rect 15 -1199 31 -1165
rect 65 -1199 81 -1165
rect 207 -1199 223 -1165
rect 257 -1199 273 -1165
rect 399 -1199 415 -1165
rect 449 -1199 465 -1165
rect -707 -1267 -673 -1205
rect 673 -1267 707 -1205
rect -707 -1301 -611 -1267
rect 611 -1301 707 -1267
<< viali >>
rect -545 1165 -511 1199
rect -353 1165 -319 1199
rect -161 1165 -127 1199
rect 31 1165 65 1199
rect 223 1165 257 1199
rect 415 1165 449 1199
rect -593 739 -559 1115
rect -497 739 -463 1115
rect -401 739 -367 1115
rect -305 739 -271 1115
rect -209 739 -175 1115
rect -113 739 -79 1115
rect -17 739 17 1115
rect 79 739 113 1115
rect 175 739 209 1115
rect 271 739 305 1115
rect 367 739 401 1115
rect 463 739 497 1115
rect 559 739 593 1115
rect -449 655 -415 689
rect -257 655 -223 689
rect -65 655 -31 689
rect 127 655 161 689
rect 319 655 353 689
rect 511 655 545 689
rect -449 547 -415 581
rect -257 547 -223 581
rect -65 547 -31 581
rect 127 547 161 581
rect 319 547 353 581
rect 511 547 545 581
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect -449 -581 -415 -547
rect -257 -581 -223 -547
rect -65 -581 -31 -547
rect 127 -581 161 -547
rect 319 -581 353 -547
rect 511 -581 545 -547
rect -449 -689 -415 -655
rect -257 -689 -223 -655
rect -65 -689 -31 -655
rect 127 -689 161 -655
rect 319 -689 353 -655
rect 511 -689 545 -655
rect -593 -1115 -559 -739
rect -497 -1115 -463 -739
rect -401 -1115 -367 -739
rect -305 -1115 -271 -739
rect -209 -1115 -175 -739
rect -113 -1115 -79 -739
rect -17 -1115 17 -739
rect 79 -1115 113 -739
rect 175 -1115 209 -739
rect 271 -1115 305 -739
rect 367 -1115 401 -739
rect 463 -1115 497 -739
rect 559 -1115 593 -739
rect -545 -1199 -511 -1165
rect -353 -1199 -319 -1165
rect -161 -1199 -127 -1165
rect 31 -1199 65 -1165
rect 223 -1199 257 -1165
rect 415 -1199 449 -1165
<< metal1 >>
rect -557 1199 -499 1205
rect -557 1165 -545 1199
rect -511 1165 -499 1199
rect -557 1159 -499 1165
rect -365 1199 -307 1205
rect -365 1165 -353 1199
rect -319 1165 -307 1199
rect -365 1159 -307 1165
rect -173 1199 -115 1205
rect -173 1165 -161 1199
rect -127 1165 -115 1199
rect -173 1159 -115 1165
rect 19 1199 77 1205
rect 19 1165 31 1199
rect 65 1165 77 1199
rect 19 1159 77 1165
rect 211 1199 269 1205
rect 211 1165 223 1199
rect 257 1165 269 1199
rect 211 1159 269 1165
rect 403 1199 461 1205
rect 403 1165 415 1199
rect 449 1165 461 1199
rect 403 1159 461 1165
rect -599 1115 -553 1127
rect -599 739 -593 1115
rect -559 739 -553 1115
rect -599 727 -553 739
rect -503 1115 -457 1127
rect -503 739 -497 1115
rect -463 739 -457 1115
rect -503 727 -457 739
rect -407 1115 -361 1127
rect -407 739 -401 1115
rect -367 739 -361 1115
rect -407 727 -361 739
rect -311 1115 -265 1127
rect -311 739 -305 1115
rect -271 739 -265 1115
rect -311 727 -265 739
rect -215 1115 -169 1127
rect -215 739 -209 1115
rect -175 739 -169 1115
rect -215 727 -169 739
rect -119 1115 -73 1127
rect -119 739 -113 1115
rect -79 739 -73 1115
rect -119 727 -73 739
rect -23 1115 23 1127
rect -23 739 -17 1115
rect 17 739 23 1115
rect -23 727 23 739
rect 73 1115 119 1127
rect 73 739 79 1115
rect 113 739 119 1115
rect 73 727 119 739
rect 169 1115 215 1127
rect 169 739 175 1115
rect 209 739 215 1115
rect 169 727 215 739
rect 265 1115 311 1127
rect 265 739 271 1115
rect 305 739 311 1115
rect 265 727 311 739
rect 361 1115 407 1127
rect 361 739 367 1115
rect 401 739 407 1115
rect 361 727 407 739
rect 457 1115 503 1127
rect 457 739 463 1115
rect 497 739 503 1115
rect 457 727 503 739
rect 553 1115 599 1127
rect 553 739 559 1115
rect 593 739 599 1115
rect 553 727 599 739
rect -461 689 -403 695
rect -461 655 -449 689
rect -415 655 -403 689
rect -461 649 -403 655
rect -269 689 -211 695
rect -269 655 -257 689
rect -223 655 -211 689
rect -269 649 -211 655
rect -77 689 -19 695
rect -77 655 -65 689
rect -31 655 -19 689
rect -77 649 -19 655
rect 115 689 173 695
rect 115 655 127 689
rect 161 655 173 689
rect 115 649 173 655
rect 307 689 365 695
rect 307 655 319 689
rect 353 655 365 689
rect 307 649 365 655
rect 499 689 557 695
rect 499 655 511 689
rect 545 655 557 689
rect 499 649 557 655
rect -461 581 -403 587
rect -461 547 -449 581
rect -415 547 -403 581
rect -461 541 -403 547
rect -269 581 -211 587
rect -269 547 -257 581
rect -223 547 -211 581
rect -269 541 -211 547
rect -77 581 -19 587
rect -77 547 -65 581
rect -31 547 -19 581
rect -77 541 -19 547
rect 115 581 173 587
rect 115 547 127 581
rect 161 547 173 581
rect 115 541 173 547
rect 307 581 365 587
rect 307 547 319 581
rect 353 547 365 581
rect 307 541 365 547
rect 499 581 557 587
rect 499 547 511 581
rect 545 547 557 581
rect 499 541 557 547
rect -599 497 -553 509
rect -599 121 -593 497
rect -559 121 -553 497
rect -599 109 -553 121
rect -503 497 -457 509
rect -503 121 -497 497
rect -463 121 -457 497
rect -503 109 -457 121
rect -407 497 -361 509
rect -407 121 -401 497
rect -367 121 -361 497
rect -407 109 -361 121
rect -311 497 -265 509
rect -311 121 -305 497
rect -271 121 -265 497
rect -311 109 -265 121
rect -215 497 -169 509
rect -215 121 -209 497
rect -175 121 -169 497
rect -215 109 -169 121
rect -119 497 -73 509
rect -119 121 -113 497
rect -79 121 -73 497
rect -119 109 -73 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 73 497 119 509
rect 73 121 79 497
rect 113 121 119 497
rect 73 109 119 121
rect 169 497 215 509
rect 169 121 175 497
rect 209 121 215 497
rect 169 109 215 121
rect 265 497 311 509
rect 265 121 271 497
rect 305 121 311 497
rect 265 109 311 121
rect 361 497 407 509
rect 361 121 367 497
rect 401 121 407 497
rect 361 109 407 121
rect 457 497 503 509
rect 457 121 463 497
rect 497 121 503 497
rect 457 109 503 121
rect 553 497 599 509
rect 553 121 559 497
rect 593 121 599 497
rect 553 109 599 121
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect -599 -121 -553 -109
rect -599 -497 -593 -121
rect -559 -497 -553 -121
rect -599 -509 -553 -497
rect -503 -121 -457 -109
rect -503 -497 -497 -121
rect -463 -497 -457 -121
rect -503 -509 -457 -497
rect -407 -121 -361 -109
rect -407 -497 -401 -121
rect -367 -497 -361 -121
rect -407 -509 -361 -497
rect -311 -121 -265 -109
rect -311 -497 -305 -121
rect -271 -497 -265 -121
rect -311 -509 -265 -497
rect -215 -121 -169 -109
rect -215 -497 -209 -121
rect -175 -497 -169 -121
rect -215 -509 -169 -497
rect -119 -121 -73 -109
rect -119 -497 -113 -121
rect -79 -497 -73 -121
rect -119 -509 -73 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 73 -121 119 -109
rect 73 -497 79 -121
rect 113 -497 119 -121
rect 73 -509 119 -497
rect 169 -121 215 -109
rect 169 -497 175 -121
rect 209 -497 215 -121
rect 169 -509 215 -497
rect 265 -121 311 -109
rect 265 -497 271 -121
rect 305 -497 311 -121
rect 265 -509 311 -497
rect 361 -121 407 -109
rect 361 -497 367 -121
rect 401 -497 407 -121
rect 361 -509 407 -497
rect 457 -121 503 -109
rect 457 -497 463 -121
rect 497 -497 503 -121
rect 457 -509 503 -497
rect 553 -121 599 -109
rect 553 -497 559 -121
rect 593 -497 599 -121
rect 553 -509 599 -497
rect -461 -547 -403 -541
rect -461 -581 -449 -547
rect -415 -581 -403 -547
rect -461 -587 -403 -581
rect -269 -547 -211 -541
rect -269 -581 -257 -547
rect -223 -581 -211 -547
rect -269 -587 -211 -581
rect -77 -547 -19 -541
rect -77 -581 -65 -547
rect -31 -581 -19 -547
rect -77 -587 -19 -581
rect 115 -547 173 -541
rect 115 -581 127 -547
rect 161 -581 173 -547
rect 115 -587 173 -581
rect 307 -547 365 -541
rect 307 -581 319 -547
rect 353 -581 365 -547
rect 307 -587 365 -581
rect 499 -547 557 -541
rect 499 -581 511 -547
rect 545 -581 557 -547
rect 499 -587 557 -581
rect -461 -655 -403 -649
rect -461 -689 -449 -655
rect -415 -689 -403 -655
rect -461 -695 -403 -689
rect -269 -655 -211 -649
rect -269 -689 -257 -655
rect -223 -689 -211 -655
rect -269 -695 -211 -689
rect -77 -655 -19 -649
rect -77 -689 -65 -655
rect -31 -689 -19 -655
rect -77 -695 -19 -689
rect 115 -655 173 -649
rect 115 -689 127 -655
rect 161 -689 173 -655
rect 115 -695 173 -689
rect 307 -655 365 -649
rect 307 -689 319 -655
rect 353 -689 365 -655
rect 307 -695 365 -689
rect 499 -655 557 -649
rect 499 -689 511 -655
rect 545 -689 557 -655
rect 499 -695 557 -689
rect -599 -739 -553 -727
rect -599 -1115 -593 -739
rect -559 -1115 -553 -739
rect -599 -1127 -553 -1115
rect -503 -739 -457 -727
rect -503 -1115 -497 -739
rect -463 -1115 -457 -739
rect -503 -1127 -457 -1115
rect -407 -739 -361 -727
rect -407 -1115 -401 -739
rect -367 -1115 -361 -739
rect -407 -1127 -361 -1115
rect -311 -739 -265 -727
rect -311 -1115 -305 -739
rect -271 -1115 -265 -739
rect -311 -1127 -265 -1115
rect -215 -739 -169 -727
rect -215 -1115 -209 -739
rect -175 -1115 -169 -739
rect -215 -1127 -169 -1115
rect -119 -739 -73 -727
rect -119 -1115 -113 -739
rect -79 -1115 -73 -739
rect -119 -1127 -73 -1115
rect -23 -739 23 -727
rect -23 -1115 -17 -739
rect 17 -1115 23 -739
rect -23 -1127 23 -1115
rect 73 -739 119 -727
rect 73 -1115 79 -739
rect 113 -1115 119 -739
rect 73 -1127 119 -1115
rect 169 -739 215 -727
rect 169 -1115 175 -739
rect 209 -1115 215 -739
rect 169 -1127 215 -1115
rect 265 -739 311 -727
rect 265 -1115 271 -739
rect 305 -1115 311 -739
rect 265 -1127 311 -1115
rect 361 -739 407 -727
rect 361 -1115 367 -739
rect 401 -1115 407 -739
rect 361 -1127 407 -1115
rect 457 -739 503 -727
rect 457 -1115 463 -739
rect 497 -1115 503 -739
rect 457 -1127 503 -1115
rect 553 -739 599 -727
rect 553 -1115 559 -739
rect 593 -1115 599 -739
rect 553 -1127 599 -1115
rect -557 -1165 -499 -1159
rect -557 -1199 -545 -1165
rect -511 -1199 -499 -1165
rect -557 -1205 -499 -1199
rect -365 -1165 -307 -1159
rect -365 -1199 -353 -1165
rect -319 -1199 -307 -1165
rect -365 -1205 -307 -1199
rect -173 -1165 -115 -1159
rect -173 -1199 -161 -1165
rect -127 -1199 -115 -1165
rect -173 -1205 -115 -1199
rect 19 -1165 77 -1159
rect 19 -1199 31 -1165
rect 65 -1199 77 -1165
rect 19 -1205 77 -1199
rect 211 -1165 269 -1159
rect 211 -1199 223 -1165
rect 257 -1199 269 -1165
rect 211 -1205 269 -1199
rect 403 -1165 461 -1159
rect 403 -1199 415 -1165
rect 449 -1199 461 -1165
rect 403 -1205 461 -1199
<< properties >>
string FIXED_BBOX -690 -1284 690 1284
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 4 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
