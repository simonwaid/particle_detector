magic
tech sky130B
magscale 1 2
timestamp 1654697436
<< pwell >>
rect -483 -410 483 410
<< nmos >>
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
<< ndiff >>
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
<< ndiffc >>
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
<< psubdiff >>
rect -447 340 -351 374
rect 351 340 447 374
rect -447 278 -413 340
rect 413 278 447 340
rect -447 -340 -413 -278
rect 413 -340 447 -278
rect -447 -374 -351 -340
rect 351 -374 447 -340
<< psubdiffcont >>
rect -351 340 351 374
rect -447 -278 -413 278
rect 413 -278 447 278
rect -351 -374 351 -340
<< poly >>
rect -287 272 -187 288
rect -287 238 -271 272
rect -203 238 -187 272
rect -287 200 -187 238
rect -129 272 -29 288
rect -129 238 -113 272
rect -45 238 -29 272
rect -129 200 -29 238
rect 29 272 129 288
rect 29 238 45 272
rect 113 238 129 272
rect 29 200 129 238
rect 187 272 287 288
rect 187 238 203 272
rect 271 238 287 272
rect 187 200 287 238
rect -287 -238 -187 -200
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -287 -288 -187 -272
rect -129 -238 -29 -200
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect -129 -288 -29 -272
rect 29 -238 129 -200
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 29 -288 129 -272
rect 187 -238 287 -200
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 187 -288 287 -272
<< polycont >>
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
<< locali >>
rect -447 340 -351 374
rect 351 340 447 374
rect -447 278 -413 340
rect 413 278 447 340
rect -287 238 -271 272
rect -203 238 -187 272
rect -129 238 -113 272
rect -45 238 -29 272
rect 29 238 45 272
rect 113 238 129 272
rect 187 238 203 272
rect 271 238 287 272
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 187 -272 203 -238
rect 271 -272 287 -238
rect -447 -340 -413 -278
rect 413 -340 447 -278
rect -447 -374 -351 -340
rect 351 -374 447 -340
<< viali >>
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
<< metal1 >>
rect -283 272 -191 278
rect -283 238 -271 272
rect -203 238 -191 272
rect -283 232 -191 238
rect -125 272 -33 278
rect -125 238 -113 272
rect -45 238 -33 272
rect -125 232 -33 238
rect 33 272 125 278
rect 33 238 45 272
rect 113 238 125 272
rect 33 232 125 238
rect 191 272 283 278
rect 191 238 203 272
rect 271 238 283 272
rect 191 232 283 238
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect -283 -238 -191 -232
rect -283 -272 -271 -238
rect -203 -272 -191 -238
rect -283 -278 -191 -272
rect -125 -238 -33 -232
rect -125 -272 -113 -238
rect -45 -272 -33 -238
rect -125 -278 -33 -272
rect 33 -238 125 -232
rect 33 -272 45 -238
rect 113 -272 125 -238
rect 33 -278 125 -272
rect 191 -238 283 -232
rect 191 -272 203 -238
rect 271 -272 283 -238
rect 191 -278 283 -272
<< properties >>
string FIXED_BBOX -430 -357 430 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
