magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< error_p >>
rect -479 281 -417 287
rect -351 281 -289 287
rect -223 281 -161 287
rect -95 281 -33 287
rect 33 281 95 287
rect 161 281 223 287
rect 289 281 351 287
rect 417 281 479 287
rect -479 247 -467 281
rect -351 247 -339 281
rect -223 247 -211 281
rect -95 247 -83 281
rect 33 247 45 281
rect 161 247 173 281
rect 289 247 301 281
rect 417 247 429 281
rect -479 241 -417 247
rect -351 241 -289 247
rect -223 241 -161 247
rect -95 241 -33 247
rect 33 241 95 247
rect 161 241 223 247
rect 289 241 351 247
rect 417 241 479 247
rect -479 -247 -417 -241
rect -351 -247 -289 -241
rect -223 -247 -161 -241
rect -95 -247 -33 -241
rect 33 -247 95 -241
rect 161 -247 223 -241
rect 289 -247 351 -241
rect 417 -247 479 -241
rect -479 -281 -467 -247
rect -351 -281 -339 -247
rect -223 -281 -211 -247
rect -95 -281 -83 -247
rect 33 -281 45 -247
rect 161 -281 173 -247
rect 289 -281 301 -247
rect 417 -281 429 -247
rect -479 -287 -417 -281
rect -351 -287 -289 -281
rect -223 -287 -161 -281
rect -95 -287 -33 -281
rect 33 -287 95 -281
rect 161 -287 223 -281
rect 289 -287 351 -281
rect 417 -287 479 -281
<< nwell >>
rect -679 -419 679 419
<< pmoslvt >>
rect -483 -200 -413 200
rect -355 -200 -285 200
rect -227 -200 -157 200
rect -99 -200 -29 200
rect 29 -200 99 200
rect 157 -200 227 200
rect 285 -200 355 200
rect 413 -200 483 200
<< pdiff >>
rect -541 188 -483 200
rect -541 -188 -529 188
rect -495 -188 -483 188
rect -541 -200 -483 -188
rect -413 188 -355 200
rect -413 -188 -401 188
rect -367 -188 -355 188
rect -413 -200 -355 -188
rect -285 188 -227 200
rect -285 -188 -273 188
rect -239 -188 -227 188
rect -285 -200 -227 -188
rect -157 188 -99 200
rect -157 -188 -145 188
rect -111 -188 -99 188
rect -157 -200 -99 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 99 188 157 200
rect 99 -188 111 188
rect 145 -188 157 188
rect 99 -200 157 -188
rect 227 188 285 200
rect 227 -188 239 188
rect 273 -188 285 188
rect 227 -200 285 -188
rect 355 188 413 200
rect 355 -188 367 188
rect 401 -188 413 188
rect 355 -200 413 -188
rect 483 188 541 200
rect 483 -188 495 188
rect 529 -188 541 188
rect 483 -200 541 -188
<< pdiffc >>
rect -529 -188 -495 188
rect -401 -188 -367 188
rect -273 -188 -239 188
rect -145 -188 -111 188
rect -17 -188 17 188
rect 111 -188 145 188
rect 239 -188 273 188
rect 367 -188 401 188
rect 495 -188 529 188
<< nsubdiff >>
rect -643 349 -547 383
rect 547 349 643 383
rect -643 287 -609 349
rect 609 287 643 349
rect -643 -349 -609 -287
rect 609 -349 643 -287
rect -643 -383 -547 -349
rect 547 -383 643 -349
<< nsubdiffcont >>
rect -547 349 547 383
rect -643 -287 -609 287
rect 609 -287 643 287
rect -547 -383 547 -349
<< poly >>
rect -483 281 -413 297
rect -483 247 -467 281
rect -429 247 -413 281
rect -483 200 -413 247
rect -355 281 -285 297
rect -355 247 -339 281
rect -301 247 -285 281
rect -355 200 -285 247
rect -227 281 -157 297
rect -227 247 -211 281
rect -173 247 -157 281
rect -227 200 -157 247
rect -99 281 -29 297
rect -99 247 -83 281
rect -45 247 -29 281
rect -99 200 -29 247
rect 29 281 99 297
rect 29 247 45 281
rect 83 247 99 281
rect 29 200 99 247
rect 157 281 227 297
rect 157 247 173 281
rect 211 247 227 281
rect 157 200 227 247
rect 285 281 355 297
rect 285 247 301 281
rect 339 247 355 281
rect 285 200 355 247
rect 413 281 483 297
rect 413 247 429 281
rect 467 247 483 281
rect 413 200 483 247
rect -483 -247 -413 -200
rect -483 -281 -467 -247
rect -429 -281 -413 -247
rect -483 -297 -413 -281
rect -355 -247 -285 -200
rect -355 -281 -339 -247
rect -301 -281 -285 -247
rect -355 -297 -285 -281
rect -227 -247 -157 -200
rect -227 -281 -211 -247
rect -173 -281 -157 -247
rect -227 -297 -157 -281
rect -99 -247 -29 -200
rect -99 -281 -83 -247
rect -45 -281 -29 -247
rect -99 -297 -29 -281
rect 29 -247 99 -200
rect 29 -281 45 -247
rect 83 -281 99 -247
rect 29 -297 99 -281
rect 157 -247 227 -200
rect 157 -281 173 -247
rect 211 -281 227 -247
rect 157 -297 227 -281
rect 285 -247 355 -200
rect 285 -281 301 -247
rect 339 -281 355 -247
rect 285 -297 355 -281
rect 413 -247 483 -200
rect 413 -281 429 -247
rect 467 -281 483 -247
rect 413 -297 483 -281
<< polycont >>
rect -467 247 -429 281
rect -339 247 -301 281
rect -211 247 -173 281
rect -83 247 -45 281
rect 45 247 83 281
rect 173 247 211 281
rect 301 247 339 281
rect 429 247 467 281
rect -467 -281 -429 -247
rect -339 -281 -301 -247
rect -211 -281 -173 -247
rect -83 -281 -45 -247
rect 45 -281 83 -247
rect 173 -281 211 -247
rect 301 -281 339 -247
rect 429 -281 467 -247
<< locali >>
rect -643 349 -547 383
rect 547 349 643 383
rect -643 287 -609 349
rect 609 287 643 349
rect -483 247 -467 281
rect -429 247 -413 281
rect -355 247 -339 281
rect -301 247 -285 281
rect -227 247 -211 281
rect -173 247 -157 281
rect -99 247 -83 281
rect -45 247 -29 281
rect 29 247 45 281
rect 83 247 99 281
rect 157 247 173 281
rect 211 247 227 281
rect 285 247 301 281
rect 339 247 355 281
rect 413 247 429 281
rect 467 247 483 281
rect -529 188 -495 204
rect -529 -204 -495 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -273 188 -239 204
rect -273 -204 -239 -188
rect -145 188 -111 204
rect -145 -204 -111 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 111 188 145 204
rect 111 -204 145 -188
rect 239 188 273 204
rect 239 -204 273 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 495 188 529 204
rect 495 -204 529 -188
rect -483 -281 -467 -247
rect -429 -281 -413 -247
rect -355 -281 -339 -247
rect -301 -281 -285 -247
rect -227 -281 -211 -247
rect -173 -281 -157 -247
rect -99 -281 -83 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 83 -281 99 -247
rect 157 -281 173 -247
rect 211 -281 227 -247
rect 285 -281 301 -247
rect 339 -281 355 -247
rect 413 -281 429 -247
rect 467 -281 483 -247
rect -643 -349 -609 -287
rect 609 -349 643 -287
rect -643 -383 -547 -349
rect 547 -383 643 -349
<< viali >>
rect -467 247 -429 281
rect -339 247 -301 281
rect -211 247 -173 281
rect -83 247 -45 281
rect 45 247 83 281
rect 173 247 211 281
rect 301 247 339 281
rect 429 247 467 281
rect -529 -188 -495 188
rect -401 -188 -367 188
rect -273 -188 -239 188
rect -145 -188 -111 188
rect -17 -188 17 188
rect 111 -188 145 188
rect 239 -188 273 188
rect 367 -188 401 188
rect 495 -188 529 188
rect -467 -281 -429 -247
rect -339 -281 -301 -247
rect -211 -281 -173 -247
rect -83 -281 -45 -247
rect 45 -281 83 -247
rect 173 -281 211 -247
rect 301 -281 339 -247
rect 429 -281 467 -247
<< metal1 >>
rect -479 281 -417 287
rect -479 247 -467 281
rect -429 247 -417 281
rect -479 241 -417 247
rect -351 281 -289 287
rect -351 247 -339 281
rect -301 247 -289 281
rect -351 241 -289 247
rect -223 281 -161 287
rect -223 247 -211 281
rect -173 247 -161 281
rect -223 241 -161 247
rect -95 281 -33 287
rect -95 247 -83 281
rect -45 247 -33 281
rect -95 241 -33 247
rect 33 281 95 287
rect 33 247 45 281
rect 83 247 95 281
rect 33 241 95 247
rect 161 281 223 287
rect 161 247 173 281
rect 211 247 223 281
rect 161 241 223 247
rect 289 281 351 287
rect 289 247 301 281
rect 339 247 351 281
rect 289 241 351 247
rect 417 281 479 287
rect 417 247 429 281
rect 467 247 479 281
rect 417 241 479 247
rect -535 188 -489 200
rect -535 -188 -529 188
rect -495 -188 -489 188
rect -535 -200 -489 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -279 188 -233 200
rect -279 -188 -273 188
rect -239 -188 -233 188
rect -279 -200 -233 -188
rect -151 188 -105 200
rect -151 -188 -145 188
rect -111 -188 -105 188
rect -151 -200 -105 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 105 188 151 200
rect 105 -188 111 188
rect 145 -188 151 188
rect 105 -200 151 -188
rect 233 188 279 200
rect 233 -188 239 188
rect 273 -188 279 188
rect 233 -200 279 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 489 188 535 200
rect 489 -188 495 188
rect 529 -188 535 188
rect 489 -200 535 -188
rect -479 -247 -417 -241
rect -479 -281 -467 -247
rect -429 -281 -417 -247
rect -479 -287 -417 -281
rect -351 -247 -289 -241
rect -351 -281 -339 -247
rect -301 -281 -289 -247
rect -351 -287 -289 -281
rect -223 -247 -161 -241
rect -223 -281 -211 -247
rect -173 -281 -161 -247
rect -223 -287 -161 -281
rect -95 -247 -33 -241
rect -95 -281 -83 -247
rect -45 -281 -33 -247
rect -95 -287 -33 -281
rect 33 -247 95 -241
rect 33 -281 45 -247
rect 83 -281 95 -247
rect 33 -287 95 -281
rect 161 -247 223 -241
rect 161 -281 173 -247
rect 211 -281 223 -247
rect 161 -287 223 -281
rect 289 -247 351 -241
rect 289 -281 301 -247
rect 339 -281 351 -247
rect 289 -287 351 -281
rect 417 -247 479 -241
rect 417 -281 429 -247
rect 467 -281 479 -247
rect 417 -287 479 -281
<< properties >>
string FIXED_BBOX -626 -366 626 366
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2 l 0.35 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
