magic
tech sky130A
magscale 1 2
timestamp 1647868710
<< pwell >>
rect -1431 -2573 1431 2573
<< nmos >>
rect -1235 1963 -1135 2363
rect -1077 1963 -977 2363
rect -919 1963 -819 2363
rect -761 1963 -661 2363
rect -603 1963 -503 2363
rect -445 1963 -345 2363
rect -287 1963 -187 2363
rect -129 1963 -29 2363
rect 29 1963 129 2363
rect 187 1963 287 2363
rect 345 1963 445 2363
rect 503 1963 603 2363
rect 661 1963 761 2363
rect 819 1963 919 2363
rect 977 1963 1077 2363
rect 1135 1963 1235 2363
rect -1235 1345 -1135 1745
rect -1077 1345 -977 1745
rect -919 1345 -819 1745
rect -761 1345 -661 1745
rect -603 1345 -503 1745
rect -445 1345 -345 1745
rect -287 1345 -187 1745
rect -129 1345 -29 1745
rect 29 1345 129 1745
rect 187 1345 287 1745
rect 345 1345 445 1745
rect 503 1345 603 1745
rect 661 1345 761 1745
rect 819 1345 919 1745
rect 977 1345 1077 1745
rect 1135 1345 1235 1745
rect -1235 727 -1135 1127
rect -1077 727 -977 1127
rect -919 727 -819 1127
rect -761 727 -661 1127
rect -603 727 -503 1127
rect -445 727 -345 1127
rect -287 727 -187 1127
rect -129 727 -29 1127
rect 29 727 129 1127
rect 187 727 287 1127
rect 345 727 445 1127
rect 503 727 603 1127
rect 661 727 761 1127
rect 819 727 919 1127
rect 977 727 1077 1127
rect 1135 727 1235 1127
rect -1235 109 -1135 509
rect -1077 109 -977 509
rect -919 109 -819 509
rect -761 109 -661 509
rect -603 109 -503 509
rect -445 109 -345 509
rect -287 109 -187 509
rect -129 109 -29 509
rect 29 109 129 509
rect 187 109 287 509
rect 345 109 445 509
rect 503 109 603 509
rect 661 109 761 509
rect 819 109 919 509
rect 977 109 1077 509
rect 1135 109 1235 509
rect -1235 -509 -1135 -109
rect -1077 -509 -977 -109
rect -919 -509 -819 -109
rect -761 -509 -661 -109
rect -603 -509 -503 -109
rect -445 -509 -345 -109
rect -287 -509 -187 -109
rect -129 -509 -29 -109
rect 29 -509 129 -109
rect 187 -509 287 -109
rect 345 -509 445 -109
rect 503 -509 603 -109
rect 661 -509 761 -109
rect 819 -509 919 -109
rect 977 -509 1077 -109
rect 1135 -509 1235 -109
rect -1235 -1127 -1135 -727
rect -1077 -1127 -977 -727
rect -919 -1127 -819 -727
rect -761 -1127 -661 -727
rect -603 -1127 -503 -727
rect -445 -1127 -345 -727
rect -287 -1127 -187 -727
rect -129 -1127 -29 -727
rect 29 -1127 129 -727
rect 187 -1127 287 -727
rect 345 -1127 445 -727
rect 503 -1127 603 -727
rect 661 -1127 761 -727
rect 819 -1127 919 -727
rect 977 -1127 1077 -727
rect 1135 -1127 1235 -727
rect -1235 -1745 -1135 -1345
rect -1077 -1745 -977 -1345
rect -919 -1745 -819 -1345
rect -761 -1745 -661 -1345
rect -603 -1745 -503 -1345
rect -445 -1745 -345 -1345
rect -287 -1745 -187 -1345
rect -129 -1745 -29 -1345
rect 29 -1745 129 -1345
rect 187 -1745 287 -1345
rect 345 -1745 445 -1345
rect 503 -1745 603 -1345
rect 661 -1745 761 -1345
rect 819 -1745 919 -1345
rect 977 -1745 1077 -1345
rect 1135 -1745 1235 -1345
rect -1235 -2363 -1135 -1963
rect -1077 -2363 -977 -1963
rect -919 -2363 -819 -1963
rect -761 -2363 -661 -1963
rect -603 -2363 -503 -1963
rect -445 -2363 -345 -1963
rect -287 -2363 -187 -1963
rect -129 -2363 -29 -1963
rect 29 -2363 129 -1963
rect 187 -2363 287 -1963
rect 345 -2363 445 -1963
rect 503 -2363 603 -1963
rect 661 -2363 761 -1963
rect 819 -2363 919 -1963
rect 977 -2363 1077 -1963
rect 1135 -2363 1235 -1963
<< ndiff >>
rect -1293 2351 -1235 2363
rect -1293 1975 -1281 2351
rect -1247 1975 -1235 2351
rect -1293 1963 -1235 1975
rect -1135 2351 -1077 2363
rect -1135 1975 -1123 2351
rect -1089 1975 -1077 2351
rect -1135 1963 -1077 1975
rect -977 2351 -919 2363
rect -977 1975 -965 2351
rect -931 1975 -919 2351
rect -977 1963 -919 1975
rect -819 2351 -761 2363
rect -819 1975 -807 2351
rect -773 1975 -761 2351
rect -819 1963 -761 1975
rect -661 2351 -603 2363
rect -661 1975 -649 2351
rect -615 1975 -603 2351
rect -661 1963 -603 1975
rect -503 2351 -445 2363
rect -503 1975 -491 2351
rect -457 1975 -445 2351
rect -503 1963 -445 1975
rect -345 2351 -287 2363
rect -345 1975 -333 2351
rect -299 1975 -287 2351
rect -345 1963 -287 1975
rect -187 2351 -129 2363
rect -187 1975 -175 2351
rect -141 1975 -129 2351
rect -187 1963 -129 1975
rect -29 2351 29 2363
rect -29 1975 -17 2351
rect 17 1975 29 2351
rect -29 1963 29 1975
rect 129 2351 187 2363
rect 129 1975 141 2351
rect 175 1975 187 2351
rect 129 1963 187 1975
rect 287 2351 345 2363
rect 287 1975 299 2351
rect 333 1975 345 2351
rect 287 1963 345 1975
rect 445 2351 503 2363
rect 445 1975 457 2351
rect 491 1975 503 2351
rect 445 1963 503 1975
rect 603 2351 661 2363
rect 603 1975 615 2351
rect 649 1975 661 2351
rect 603 1963 661 1975
rect 761 2351 819 2363
rect 761 1975 773 2351
rect 807 1975 819 2351
rect 761 1963 819 1975
rect 919 2351 977 2363
rect 919 1975 931 2351
rect 965 1975 977 2351
rect 919 1963 977 1975
rect 1077 2351 1135 2363
rect 1077 1975 1089 2351
rect 1123 1975 1135 2351
rect 1077 1963 1135 1975
rect 1235 2351 1293 2363
rect 1235 1975 1247 2351
rect 1281 1975 1293 2351
rect 1235 1963 1293 1975
rect -1293 1733 -1235 1745
rect -1293 1357 -1281 1733
rect -1247 1357 -1235 1733
rect -1293 1345 -1235 1357
rect -1135 1733 -1077 1745
rect -1135 1357 -1123 1733
rect -1089 1357 -1077 1733
rect -1135 1345 -1077 1357
rect -977 1733 -919 1745
rect -977 1357 -965 1733
rect -931 1357 -919 1733
rect -977 1345 -919 1357
rect -819 1733 -761 1745
rect -819 1357 -807 1733
rect -773 1357 -761 1733
rect -819 1345 -761 1357
rect -661 1733 -603 1745
rect -661 1357 -649 1733
rect -615 1357 -603 1733
rect -661 1345 -603 1357
rect -503 1733 -445 1745
rect -503 1357 -491 1733
rect -457 1357 -445 1733
rect -503 1345 -445 1357
rect -345 1733 -287 1745
rect -345 1357 -333 1733
rect -299 1357 -287 1733
rect -345 1345 -287 1357
rect -187 1733 -129 1745
rect -187 1357 -175 1733
rect -141 1357 -129 1733
rect -187 1345 -129 1357
rect -29 1733 29 1745
rect -29 1357 -17 1733
rect 17 1357 29 1733
rect -29 1345 29 1357
rect 129 1733 187 1745
rect 129 1357 141 1733
rect 175 1357 187 1733
rect 129 1345 187 1357
rect 287 1733 345 1745
rect 287 1357 299 1733
rect 333 1357 345 1733
rect 287 1345 345 1357
rect 445 1733 503 1745
rect 445 1357 457 1733
rect 491 1357 503 1733
rect 445 1345 503 1357
rect 603 1733 661 1745
rect 603 1357 615 1733
rect 649 1357 661 1733
rect 603 1345 661 1357
rect 761 1733 819 1745
rect 761 1357 773 1733
rect 807 1357 819 1733
rect 761 1345 819 1357
rect 919 1733 977 1745
rect 919 1357 931 1733
rect 965 1357 977 1733
rect 919 1345 977 1357
rect 1077 1733 1135 1745
rect 1077 1357 1089 1733
rect 1123 1357 1135 1733
rect 1077 1345 1135 1357
rect 1235 1733 1293 1745
rect 1235 1357 1247 1733
rect 1281 1357 1293 1733
rect 1235 1345 1293 1357
rect -1293 1115 -1235 1127
rect -1293 739 -1281 1115
rect -1247 739 -1235 1115
rect -1293 727 -1235 739
rect -1135 1115 -1077 1127
rect -1135 739 -1123 1115
rect -1089 739 -1077 1115
rect -1135 727 -1077 739
rect -977 1115 -919 1127
rect -977 739 -965 1115
rect -931 739 -919 1115
rect -977 727 -919 739
rect -819 1115 -761 1127
rect -819 739 -807 1115
rect -773 739 -761 1115
rect -819 727 -761 739
rect -661 1115 -603 1127
rect -661 739 -649 1115
rect -615 739 -603 1115
rect -661 727 -603 739
rect -503 1115 -445 1127
rect -503 739 -491 1115
rect -457 739 -445 1115
rect -503 727 -445 739
rect -345 1115 -287 1127
rect -345 739 -333 1115
rect -299 739 -287 1115
rect -345 727 -287 739
rect -187 1115 -129 1127
rect -187 739 -175 1115
rect -141 739 -129 1115
rect -187 727 -129 739
rect -29 1115 29 1127
rect -29 739 -17 1115
rect 17 739 29 1115
rect -29 727 29 739
rect 129 1115 187 1127
rect 129 739 141 1115
rect 175 739 187 1115
rect 129 727 187 739
rect 287 1115 345 1127
rect 287 739 299 1115
rect 333 739 345 1115
rect 287 727 345 739
rect 445 1115 503 1127
rect 445 739 457 1115
rect 491 739 503 1115
rect 445 727 503 739
rect 603 1115 661 1127
rect 603 739 615 1115
rect 649 739 661 1115
rect 603 727 661 739
rect 761 1115 819 1127
rect 761 739 773 1115
rect 807 739 819 1115
rect 761 727 819 739
rect 919 1115 977 1127
rect 919 739 931 1115
rect 965 739 977 1115
rect 919 727 977 739
rect 1077 1115 1135 1127
rect 1077 739 1089 1115
rect 1123 739 1135 1115
rect 1077 727 1135 739
rect 1235 1115 1293 1127
rect 1235 739 1247 1115
rect 1281 739 1293 1115
rect 1235 727 1293 739
rect -1293 497 -1235 509
rect -1293 121 -1281 497
rect -1247 121 -1235 497
rect -1293 109 -1235 121
rect -1135 497 -1077 509
rect -1135 121 -1123 497
rect -1089 121 -1077 497
rect -1135 109 -1077 121
rect -977 497 -919 509
rect -977 121 -965 497
rect -931 121 -919 497
rect -977 109 -919 121
rect -819 497 -761 509
rect -819 121 -807 497
rect -773 121 -761 497
rect -819 109 -761 121
rect -661 497 -603 509
rect -661 121 -649 497
rect -615 121 -603 497
rect -661 109 -603 121
rect -503 497 -445 509
rect -503 121 -491 497
rect -457 121 -445 497
rect -503 109 -445 121
rect -345 497 -287 509
rect -345 121 -333 497
rect -299 121 -287 497
rect -345 109 -287 121
rect -187 497 -129 509
rect -187 121 -175 497
rect -141 121 -129 497
rect -187 109 -129 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 129 497 187 509
rect 129 121 141 497
rect 175 121 187 497
rect 129 109 187 121
rect 287 497 345 509
rect 287 121 299 497
rect 333 121 345 497
rect 287 109 345 121
rect 445 497 503 509
rect 445 121 457 497
rect 491 121 503 497
rect 445 109 503 121
rect 603 497 661 509
rect 603 121 615 497
rect 649 121 661 497
rect 603 109 661 121
rect 761 497 819 509
rect 761 121 773 497
rect 807 121 819 497
rect 761 109 819 121
rect 919 497 977 509
rect 919 121 931 497
rect 965 121 977 497
rect 919 109 977 121
rect 1077 497 1135 509
rect 1077 121 1089 497
rect 1123 121 1135 497
rect 1077 109 1135 121
rect 1235 497 1293 509
rect 1235 121 1247 497
rect 1281 121 1293 497
rect 1235 109 1293 121
rect -1293 -121 -1235 -109
rect -1293 -497 -1281 -121
rect -1247 -497 -1235 -121
rect -1293 -509 -1235 -497
rect -1135 -121 -1077 -109
rect -1135 -497 -1123 -121
rect -1089 -497 -1077 -121
rect -1135 -509 -1077 -497
rect -977 -121 -919 -109
rect -977 -497 -965 -121
rect -931 -497 -919 -121
rect -977 -509 -919 -497
rect -819 -121 -761 -109
rect -819 -497 -807 -121
rect -773 -497 -761 -121
rect -819 -509 -761 -497
rect -661 -121 -603 -109
rect -661 -497 -649 -121
rect -615 -497 -603 -121
rect -661 -509 -603 -497
rect -503 -121 -445 -109
rect -503 -497 -491 -121
rect -457 -497 -445 -121
rect -503 -509 -445 -497
rect -345 -121 -287 -109
rect -345 -497 -333 -121
rect -299 -497 -287 -121
rect -345 -509 -287 -497
rect -187 -121 -129 -109
rect -187 -497 -175 -121
rect -141 -497 -129 -121
rect -187 -509 -129 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 129 -121 187 -109
rect 129 -497 141 -121
rect 175 -497 187 -121
rect 129 -509 187 -497
rect 287 -121 345 -109
rect 287 -497 299 -121
rect 333 -497 345 -121
rect 287 -509 345 -497
rect 445 -121 503 -109
rect 445 -497 457 -121
rect 491 -497 503 -121
rect 445 -509 503 -497
rect 603 -121 661 -109
rect 603 -497 615 -121
rect 649 -497 661 -121
rect 603 -509 661 -497
rect 761 -121 819 -109
rect 761 -497 773 -121
rect 807 -497 819 -121
rect 761 -509 819 -497
rect 919 -121 977 -109
rect 919 -497 931 -121
rect 965 -497 977 -121
rect 919 -509 977 -497
rect 1077 -121 1135 -109
rect 1077 -497 1089 -121
rect 1123 -497 1135 -121
rect 1077 -509 1135 -497
rect 1235 -121 1293 -109
rect 1235 -497 1247 -121
rect 1281 -497 1293 -121
rect 1235 -509 1293 -497
rect -1293 -739 -1235 -727
rect -1293 -1115 -1281 -739
rect -1247 -1115 -1235 -739
rect -1293 -1127 -1235 -1115
rect -1135 -739 -1077 -727
rect -1135 -1115 -1123 -739
rect -1089 -1115 -1077 -739
rect -1135 -1127 -1077 -1115
rect -977 -739 -919 -727
rect -977 -1115 -965 -739
rect -931 -1115 -919 -739
rect -977 -1127 -919 -1115
rect -819 -739 -761 -727
rect -819 -1115 -807 -739
rect -773 -1115 -761 -739
rect -819 -1127 -761 -1115
rect -661 -739 -603 -727
rect -661 -1115 -649 -739
rect -615 -1115 -603 -739
rect -661 -1127 -603 -1115
rect -503 -739 -445 -727
rect -503 -1115 -491 -739
rect -457 -1115 -445 -739
rect -503 -1127 -445 -1115
rect -345 -739 -287 -727
rect -345 -1115 -333 -739
rect -299 -1115 -287 -739
rect -345 -1127 -287 -1115
rect -187 -739 -129 -727
rect -187 -1115 -175 -739
rect -141 -1115 -129 -739
rect -187 -1127 -129 -1115
rect -29 -739 29 -727
rect -29 -1115 -17 -739
rect 17 -1115 29 -739
rect -29 -1127 29 -1115
rect 129 -739 187 -727
rect 129 -1115 141 -739
rect 175 -1115 187 -739
rect 129 -1127 187 -1115
rect 287 -739 345 -727
rect 287 -1115 299 -739
rect 333 -1115 345 -739
rect 287 -1127 345 -1115
rect 445 -739 503 -727
rect 445 -1115 457 -739
rect 491 -1115 503 -739
rect 445 -1127 503 -1115
rect 603 -739 661 -727
rect 603 -1115 615 -739
rect 649 -1115 661 -739
rect 603 -1127 661 -1115
rect 761 -739 819 -727
rect 761 -1115 773 -739
rect 807 -1115 819 -739
rect 761 -1127 819 -1115
rect 919 -739 977 -727
rect 919 -1115 931 -739
rect 965 -1115 977 -739
rect 919 -1127 977 -1115
rect 1077 -739 1135 -727
rect 1077 -1115 1089 -739
rect 1123 -1115 1135 -739
rect 1077 -1127 1135 -1115
rect 1235 -739 1293 -727
rect 1235 -1115 1247 -739
rect 1281 -1115 1293 -739
rect 1235 -1127 1293 -1115
rect -1293 -1357 -1235 -1345
rect -1293 -1733 -1281 -1357
rect -1247 -1733 -1235 -1357
rect -1293 -1745 -1235 -1733
rect -1135 -1357 -1077 -1345
rect -1135 -1733 -1123 -1357
rect -1089 -1733 -1077 -1357
rect -1135 -1745 -1077 -1733
rect -977 -1357 -919 -1345
rect -977 -1733 -965 -1357
rect -931 -1733 -919 -1357
rect -977 -1745 -919 -1733
rect -819 -1357 -761 -1345
rect -819 -1733 -807 -1357
rect -773 -1733 -761 -1357
rect -819 -1745 -761 -1733
rect -661 -1357 -603 -1345
rect -661 -1733 -649 -1357
rect -615 -1733 -603 -1357
rect -661 -1745 -603 -1733
rect -503 -1357 -445 -1345
rect -503 -1733 -491 -1357
rect -457 -1733 -445 -1357
rect -503 -1745 -445 -1733
rect -345 -1357 -287 -1345
rect -345 -1733 -333 -1357
rect -299 -1733 -287 -1357
rect -345 -1745 -287 -1733
rect -187 -1357 -129 -1345
rect -187 -1733 -175 -1357
rect -141 -1733 -129 -1357
rect -187 -1745 -129 -1733
rect -29 -1357 29 -1345
rect -29 -1733 -17 -1357
rect 17 -1733 29 -1357
rect -29 -1745 29 -1733
rect 129 -1357 187 -1345
rect 129 -1733 141 -1357
rect 175 -1733 187 -1357
rect 129 -1745 187 -1733
rect 287 -1357 345 -1345
rect 287 -1733 299 -1357
rect 333 -1733 345 -1357
rect 287 -1745 345 -1733
rect 445 -1357 503 -1345
rect 445 -1733 457 -1357
rect 491 -1733 503 -1357
rect 445 -1745 503 -1733
rect 603 -1357 661 -1345
rect 603 -1733 615 -1357
rect 649 -1733 661 -1357
rect 603 -1745 661 -1733
rect 761 -1357 819 -1345
rect 761 -1733 773 -1357
rect 807 -1733 819 -1357
rect 761 -1745 819 -1733
rect 919 -1357 977 -1345
rect 919 -1733 931 -1357
rect 965 -1733 977 -1357
rect 919 -1745 977 -1733
rect 1077 -1357 1135 -1345
rect 1077 -1733 1089 -1357
rect 1123 -1733 1135 -1357
rect 1077 -1745 1135 -1733
rect 1235 -1357 1293 -1345
rect 1235 -1733 1247 -1357
rect 1281 -1733 1293 -1357
rect 1235 -1745 1293 -1733
rect -1293 -1975 -1235 -1963
rect -1293 -2351 -1281 -1975
rect -1247 -2351 -1235 -1975
rect -1293 -2363 -1235 -2351
rect -1135 -1975 -1077 -1963
rect -1135 -2351 -1123 -1975
rect -1089 -2351 -1077 -1975
rect -1135 -2363 -1077 -2351
rect -977 -1975 -919 -1963
rect -977 -2351 -965 -1975
rect -931 -2351 -919 -1975
rect -977 -2363 -919 -2351
rect -819 -1975 -761 -1963
rect -819 -2351 -807 -1975
rect -773 -2351 -761 -1975
rect -819 -2363 -761 -2351
rect -661 -1975 -603 -1963
rect -661 -2351 -649 -1975
rect -615 -2351 -603 -1975
rect -661 -2363 -603 -2351
rect -503 -1975 -445 -1963
rect -503 -2351 -491 -1975
rect -457 -2351 -445 -1975
rect -503 -2363 -445 -2351
rect -345 -1975 -287 -1963
rect -345 -2351 -333 -1975
rect -299 -2351 -287 -1975
rect -345 -2363 -287 -2351
rect -187 -1975 -129 -1963
rect -187 -2351 -175 -1975
rect -141 -2351 -129 -1975
rect -187 -2363 -129 -2351
rect -29 -1975 29 -1963
rect -29 -2351 -17 -1975
rect 17 -2351 29 -1975
rect -29 -2363 29 -2351
rect 129 -1975 187 -1963
rect 129 -2351 141 -1975
rect 175 -2351 187 -1975
rect 129 -2363 187 -2351
rect 287 -1975 345 -1963
rect 287 -2351 299 -1975
rect 333 -2351 345 -1975
rect 287 -2363 345 -2351
rect 445 -1975 503 -1963
rect 445 -2351 457 -1975
rect 491 -2351 503 -1975
rect 445 -2363 503 -2351
rect 603 -1975 661 -1963
rect 603 -2351 615 -1975
rect 649 -2351 661 -1975
rect 603 -2363 661 -2351
rect 761 -1975 819 -1963
rect 761 -2351 773 -1975
rect 807 -2351 819 -1975
rect 761 -2363 819 -2351
rect 919 -1975 977 -1963
rect 919 -2351 931 -1975
rect 965 -2351 977 -1975
rect 919 -2363 977 -2351
rect 1077 -1975 1135 -1963
rect 1077 -2351 1089 -1975
rect 1123 -2351 1135 -1975
rect 1077 -2363 1135 -2351
rect 1235 -1975 1293 -1963
rect 1235 -2351 1247 -1975
rect 1281 -2351 1293 -1975
rect 1235 -2363 1293 -2351
<< ndiffc >>
rect -1281 1975 -1247 2351
rect -1123 1975 -1089 2351
rect -965 1975 -931 2351
rect -807 1975 -773 2351
rect -649 1975 -615 2351
rect -491 1975 -457 2351
rect -333 1975 -299 2351
rect -175 1975 -141 2351
rect -17 1975 17 2351
rect 141 1975 175 2351
rect 299 1975 333 2351
rect 457 1975 491 2351
rect 615 1975 649 2351
rect 773 1975 807 2351
rect 931 1975 965 2351
rect 1089 1975 1123 2351
rect 1247 1975 1281 2351
rect -1281 1357 -1247 1733
rect -1123 1357 -1089 1733
rect -965 1357 -931 1733
rect -807 1357 -773 1733
rect -649 1357 -615 1733
rect -491 1357 -457 1733
rect -333 1357 -299 1733
rect -175 1357 -141 1733
rect -17 1357 17 1733
rect 141 1357 175 1733
rect 299 1357 333 1733
rect 457 1357 491 1733
rect 615 1357 649 1733
rect 773 1357 807 1733
rect 931 1357 965 1733
rect 1089 1357 1123 1733
rect 1247 1357 1281 1733
rect -1281 739 -1247 1115
rect -1123 739 -1089 1115
rect -965 739 -931 1115
rect -807 739 -773 1115
rect -649 739 -615 1115
rect -491 739 -457 1115
rect -333 739 -299 1115
rect -175 739 -141 1115
rect -17 739 17 1115
rect 141 739 175 1115
rect 299 739 333 1115
rect 457 739 491 1115
rect 615 739 649 1115
rect 773 739 807 1115
rect 931 739 965 1115
rect 1089 739 1123 1115
rect 1247 739 1281 1115
rect -1281 121 -1247 497
rect -1123 121 -1089 497
rect -965 121 -931 497
rect -807 121 -773 497
rect -649 121 -615 497
rect -491 121 -457 497
rect -333 121 -299 497
rect -175 121 -141 497
rect -17 121 17 497
rect 141 121 175 497
rect 299 121 333 497
rect 457 121 491 497
rect 615 121 649 497
rect 773 121 807 497
rect 931 121 965 497
rect 1089 121 1123 497
rect 1247 121 1281 497
rect -1281 -497 -1247 -121
rect -1123 -497 -1089 -121
rect -965 -497 -931 -121
rect -807 -497 -773 -121
rect -649 -497 -615 -121
rect -491 -497 -457 -121
rect -333 -497 -299 -121
rect -175 -497 -141 -121
rect -17 -497 17 -121
rect 141 -497 175 -121
rect 299 -497 333 -121
rect 457 -497 491 -121
rect 615 -497 649 -121
rect 773 -497 807 -121
rect 931 -497 965 -121
rect 1089 -497 1123 -121
rect 1247 -497 1281 -121
rect -1281 -1115 -1247 -739
rect -1123 -1115 -1089 -739
rect -965 -1115 -931 -739
rect -807 -1115 -773 -739
rect -649 -1115 -615 -739
rect -491 -1115 -457 -739
rect -333 -1115 -299 -739
rect -175 -1115 -141 -739
rect -17 -1115 17 -739
rect 141 -1115 175 -739
rect 299 -1115 333 -739
rect 457 -1115 491 -739
rect 615 -1115 649 -739
rect 773 -1115 807 -739
rect 931 -1115 965 -739
rect 1089 -1115 1123 -739
rect 1247 -1115 1281 -739
rect -1281 -1733 -1247 -1357
rect -1123 -1733 -1089 -1357
rect -965 -1733 -931 -1357
rect -807 -1733 -773 -1357
rect -649 -1733 -615 -1357
rect -491 -1733 -457 -1357
rect -333 -1733 -299 -1357
rect -175 -1733 -141 -1357
rect -17 -1733 17 -1357
rect 141 -1733 175 -1357
rect 299 -1733 333 -1357
rect 457 -1733 491 -1357
rect 615 -1733 649 -1357
rect 773 -1733 807 -1357
rect 931 -1733 965 -1357
rect 1089 -1733 1123 -1357
rect 1247 -1733 1281 -1357
rect -1281 -2351 -1247 -1975
rect -1123 -2351 -1089 -1975
rect -965 -2351 -931 -1975
rect -807 -2351 -773 -1975
rect -649 -2351 -615 -1975
rect -491 -2351 -457 -1975
rect -333 -2351 -299 -1975
rect -175 -2351 -141 -1975
rect -17 -2351 17 -1975
rect 141 -2351 175 -1975
rect 299 -2351 333 -1975
rect 457 -2351 491 -1975
rect 615 -2351 649 -1975
rect 773 -2351 807 -1975
rect 931 -2351 965 -1975
rect 1089 -2351 1123 -1975
rect 1247 -2351 1281 -1975
<< psubdiff >>
rect -1395 2503 -1299 2537
rect 1299 2503 1395 2537
rect -1395 2441 -1361 2503
rect 1361 2441 1395 2503
rect -1395 -2503 -1361 -2441
rect 1361 -2503 1395 -2441
rect -1395 -2537 -1299 -2503
rect 1299 -2537 1395 -2503
<< psubdiffcont >>
rect -1299 2503 1299 2537
rect -1395 -2441 -1361 2441
rect 1361 -2441 1395 2441
rect -1299 -2537 1299 -2503
<< poly >>
rect -1235 2435 -1135 2451
rect -1235 2401 -1219 2435
rect -1151 2401 -1135 2435
rect -1235 2363 -1135 2401
rect -1077 2435 -977 2451
rect -1077 2401 -1061 2435
rect -993 2401 -977 2435
rect -1077 2363 -977 2401
rect -919 2435 -819 2451
rect -919 2401 -903 2435
rect -835 2401 -819 2435
rect -919 2363 -819 2401
rect -761 2435 -661 2451
rect -761 2401 -745 2435
rect -677 2401 -661 2435
rect -761 2363 -661 2401
rect -603 2435 -503 2451
rect -603 2401 -587 2435
rect -519 2401 -503 2435
rect -603 2363 -503 2401
rect -445 2435 -345 2451
rect -445 2401 -429 2435
rect -361 2401 -345 2435
rect -445 2363 -345 2401
rect -287 2435 -187 2451
rect -287 2401 -271 2435
rect -203 2401 -187 2435
rect -287 2363 -187 2401
rect -129 2435 -29 2451
rect -129 2401 -113 2435
rect -45 2401 -29 2435
rect -129 2363 -29 2401
rect 29 2435 129 2451
rect 29 2401 45 2435
rect 113 2401 129 2435
rect 29 2363 129 2401
rect 187 2435 287 2451
rect 187 2401 203 2435
rect 271 2401 287 2435
rect 187 2363 287 2401
rect 345 2435 445 2451
rect 345 2401 361 2435
rect 429 2401 445 2435
rect 345 2363 445 2401
rect 503 2435 603 2451
rect 503 2401 519 2435
rect 587 2401 603 2435
rect 503 2363 603 2401
rect 661 2435 761 2451
rect 661 2401 677 2435
rect 745 2401 761 2435
rect 661 2363 761 2401
rect 819 2435 919 2451
rect 819 2401 835 2435
rect 903 2401 919 2435
rect 819 2363 919 2401
rect 977 2435 1077 2451
rect 977 2401 993 2435
rect 1061 2401 1077 2435
rect 977 2363 1077 2401
rect 1135 2435 1235 2451
rect 1135 2401 1151 2435
rect 1219 2401 1235 2435
rect 1135 2363 1235 2401
rect -1235 1925 -1135 1963
rect -1235 1891 -1219 1925
rect -1151 1891 -1135 1925
rect -1235 1875 -1135 1891
rect -1077 1925 -977 1963
rect -1077 1891 -1061 1925
rect -993 1891 -977 1925
rect -1077 1875 -977 1891
rect -919 1925 -819 1963
rect -919 1891 -903 1925
rect -835 1891 -819 1925
rect -919 1875 -819 1891
rect -761 1925 -661 1963
rect -761 1891 -745 1925
rect -677 1891 -661 1925
rect -761 1875 -661 1891
rect -603 1925 -503 1963
rect -603 1891 -587 1925
rect -519 1891 -503 1925
rect -603 1875 -503 1891
rect -445 1925 -345 1963
rect -445 1891 -429 1925
rect -361 1891 -345 1925
rect -445 1875 -345 1891
rect -287 1925 -187 1963
rect -287 1891 -271 1925
rect -203 1891 -187 1925
rect -287 1875 -187 1891
rect -129 1925 -29 1963
rect -129 1891 -113 1925
rect -45 1891 -29 1925
rect -129 1875 -29 1891
rect 29 1925 129 1963
rect 29 1891 45 1925
rect 113 1891 129 1925
rect 29 1875 129 1891
rect 187 1925 287 1963
rect 187 1891 203 1925
rect 271 1891 287 1925
rect 187 1875 287 1891
rect 345 1925 445 1963
rect 345 1891 361 1925
rect 429 1891 445 1925
rect 345 1875 445 1891
rect 503 1925 603 1963
rect 503 1891 519 1925
rect 587 1891 603 1925
rect 503 1875 603 1891
rect 661 1925 761 1963
rect 661 1891 677 1925
rect 745 1891 761 1925
rect 661 1875 761 1891
rect 819 1925 919 1963
rect 819 1891 835 1925
rect 903 1891 919 1925
rect 819 1875 919 1891
rect 977 1925 1077 1963
rect 977 1891 993 1925
rect 1061 1891 1077 1925
rect 977 1875 1077 1891
rect 1135 1925 1235 1963
rect 1135 1891 1151 1925
rect 1219 1891 1235 1925
rect 1135 1875 1235 1891
rect -1235 1817 -1135 1833
rect -1235 1783 -1219 1817
rect -1151 1783 -1135 1817
rect -1235 1745 -1135 1783
rect -1077 1817 -977 1833
rect -1077 1783 -1061 1817
rect -993 1783 -977 1817
rect -1077 1745 -977 1783
rect -919 1817 -819 1833
rect -919 1783 -903 1817
rect -835 1783 -819 1817
rect -919 1745 -819 1783
rect -761 1817 -661 1833
rect -761 1783 -745 1817
rect -677 1783 -661 1817
rect -761 1745 -661 1783
rect -603 1817 -503 1833
rect -603 1783 -587 1817
rect -519 1783 -503 1817
rect -603 1745 -503 1783
rect -445 1817 -345 1833
rect -445 1783 -429 1817
rect -361 1783 -345 1817
rect -445 1745 -345 1783
rect -287 1817 -187 1833
rect -287 1783 -271 1817
rect -203 1783 -187 1817
rect -287 1745 -187 1783
rect -129 1817 -29 1833
rect -129 1783 -113 1817
rect -45 1783 -29 1817
rect -129 1745 -29 1783
rect 29 1817 129 1833
rect 29 1783 45 1817
rect 113 1783 129 1817
rect 29 1745 129 1783
rect 187 1817 287 1833
rect 187 1783 203 1817
rect 271 1783 287 1817
rect 187 1745 287 1783
rect 345 1817 445 1833
rect 345 1783 361 1817
rect 429 1783 445 1817
rect 345 1745 445 1783
rect 503 1817 603 1833
rect 503 1783 519 1817
rect 587 1783 603 1817
rect 503 1745 603 1783
rect 661 1817 761 1833
rect 661 1783 677 1817
rect 745 1783 761 1817
rect 661 1745 761 1783
rect 819 1817 919 1833
rect 819 1783 835 1817
rect 903 1783 919 1817
rect 819 1745 919 1783
rect 977 1817 1077 1833
rect 977 1783 993 1817
rect 1061 1783 1077 1817
rect 977 1745 1077 1783
rect 1135 1817 1235 1833
rect 1135 1783 1151 1817
rect 1219 1783 1235 1817
rect 1135 1745 1235 1783
rect -1235 1307 -1135 1345
rect -1235 1273 -1219 1307
rect -1151 1273 -1135 1307
rect -1235 1257 -1135 1273
rect -1077 1307 -977 1345
rect -1077 1273 -1061 1307
rect -993 1273 -977 1307
rect -1077 1257 -977 1273
rect -919 1307 -819 1345
rect -919 1273 -903 1307
rect -835 1273 -819 1307
rect -919 1257 -819 1273
rect -761 1307 -661 1345
rect -761 1273 -745 1307
rect -677 1273 -661 1307
rect -761 1257 -661 1273
rect -603 1307 -503 1345
rect -603 1273 -587 1307
rect -519 1273 -503 1307
rect -603 1257 -503 1273
rect -445 1307 -345 1345
rect -445 1273 -429 1307
rect -361 1273 -345 1307
rect -445 1257 -345 1273
rect -287 1307 -187 1345
rect -287 1273 -271 1307
rect -203 1273 -187 1307
rect -287 1257 -187 1273
rect -129 1307 -29 1345
rect -129 1273 -113 1307
rect -45 1273 -29 1307
rect -129 1257 -29 1273
rect 29 1307 129 1345
rect 29 1273 45 1307
rect 113 1273 129 1307
rect 29 1257 129 1273
rect 187 1307 287 1345
rect 187 1273 203 1307
rect 271 1273 287 1307
rect 187 1257 287 1273
rect 345 1307 445 1345
rect 345 1273 361 1307
rect 429 1273 445 1307
rect 345 1257 445 1273
rect 503 1307 603 1345
rect 503 1273 519 1307
rect 587 1273 603 1307
rect 503 1257 603 1273
rect 661 1307 761 1345
rect 661 1273 677 1307
rect 745 1273 761 1307
rect 661 1257 761 1273
rect 819 1307 919 1345
rect 819 1273 835 1307
rect 903 1273 919 1307
rect 819 1257 919 1273
rect 977 1307 1077 1345
rect 977 1273 993 1307
rect 1061 1273 1077 1307
rect 977 1257 1077 1273
rect 1135 1307 1235 1345
rect 1135 1273 1151 1307
rect 1219 1273 1235 1307
rect 1135 1257 1235 1273
rect -1235 1199 -1135 1215
rect -1235 1165 -1219 1199
rect -1151 1165 -1135 1199
rect -1235 1127 -1135 1165
rect -1077 1199 -977 1215
rect -1077 1165 -1061 1199
rect -993 1165 -977 1199
rect -1077 1127 -977 1165
rect -919 1199 -819 1215
rect -919 1165 -903 1199
rect -835 1165 -819 1199
rect -919 1127 -819 1165
rect -761 1199 -661 1215
rect -761 1165 -745 1199
rect -677 1165 -661 1199
rect -761 1127 -661 1165
rect -603 1199 -503 1215
rect -603 1165 -587 1199
rect -519 1165 -503 1199
rect -603 1127 -503 1165
rect -445 1199 -345 1215
rect -445 1165 -429 1199
rect -361 1165 -345 1199
rect -445 1127 -345 1165
rect -287 1199 -187 1215
rect -287 1165 -271 1199
rect -203 1165 -187 1199
rect -287 1127 -187 1165
rect -129 1199 -29 1215
rect -129 1165 -113 1199
rect -45 1165 -29 1199
rect -129 1127 -29 1165
rect 29 1199 129 1215
rect 29 1165 45 1199
rect 113 1165 129 1199
rect 29 1127 129 1165
rect 187 1199 287 1215
rect 187 1165 203 1199
rect 271 1165 287 1199
rect 187 1127 287 1165
rect 345 1199 445 1215
rect 345 1165 361 1199
rect 429 1165 445 1199
rect 345 1127 445 1165
rect 503 1199 603 1215
rect 503 1165 519 1199
rect 587 1165 603 1199
rect 503 1127 603 1165
rect 661 1199 761 1215
rect 661 1165 677 1199
rect 745 1165 761 1199
rect 661 1127 761 1165
rect 819 1199 919 1215
rect 819 1165 835 1199
rect 903 1165 919 1199
rect 819 1127 919 1165
rect 977 1199 1077 1215
rect 977 1165 993 1199
rect 1061 1165 1077 1199
rect 977 1127 1077 1165
rect 1135 1199 1235 1215
rect 1135 1165 1151 1199
rect 1219 1165 1235 1199
rect 1135 1127 1235 1165
rect -1235 689 -1135 727
rect -1235 655 -1219 689
rect -1151 655 -1135 689
rect -1235 639 -1135 655
rect -1077 689 -977 727
rect -1077 655 -1061 689
rect -993 655 -977 689
rect -1077 639 -977 655
rect -919 689 -819 727
rect -919 655 -903 689
rect -835 655 -819 689
rect -919 639 -819 655
rect -761 689 -661 727
rect -761 655 -745 689
rect -677 655 -661 689
rect -761 639 -661 655
rect -603 689 -503 727
rect -603 655 -587 689
rect -519 655 -503 689
rect -603 639 -503 655
rect -445 689 -345 727
rect -445 655 -429 689
rect -361 655 -345 689
rect -445 639 -345 655
rect -287 689 -187 727
rect -287 655 -271 689
rect -203 655 -187 689
rect -287 639 -187 655
rect -129 689 -29 727
rect -129 655 -113 689
rect -45 655 -29 689
rect -129 639 -29 655
rect 29 689 129 727
rect 29 655 45 689
rect 113 655 129 689
rect 29 639 129 655
rect 187 689 287 727
rect 187 655 203 689
rect 271 655 287 689
rect 187 639 287 655
rect 345 689 445 727
rect 345 655 361 689
rect 429 655 445 689
rect 345 639 445 655
rect 503 689 603 727
rect 503 655 519 689
rect 587 655 603 689
rect 503 639 603 655
rect 661 689 761 727
rect 661 655 677 689
rect 745 655 761 689
rect 661 639 761 655
rect 819 689 919 727
rect 819 655 835 689
rect 903 655 919 689
rect 819 639 919 655
rect 977 689 1077 727
rect 977 655 993 689
rect 1061 655 1077 689
rect 977 639 1077 655
rect 1135 689 1235 727
rect 1135 655 1151 689
rect 1219 655 1235 689
rect 1135 639 1235 655
rect -1235 581 -1135 597
rect -1235 547 -1219 581
rect -1151 547 -1135 581
rect -1235 509 -1135 547
rect -1077 581 -977 597
rect -1077 547 -1061 581
rect -993 547 -977 581
rect -1077 509 -977 547
rect -919 581 -819 597
rect -919 547 -903 581
rect -835 547 -819 581
rect -919 509 -819 547
rect -761 581 -661 597
rect -761 547 -745 581
rect -677 547 -661 581
rect -761 509 -661 547
rect -603 581 -503 597
rect -603 547 -587 581
rect -519 547 -503 581
rect -603 509 -503 547
rect -445 581 -345 597
rect -445 547 -429 581
rect -361 547 -345 581
rect -445 509 -345 547
rect -287 581 -187 597
rect -287 547 -271 581
rect -203 547 -187 581
rect -287 509 -187 547
rect -129 581 -29 597
rect -129 547 -113 581
rect -45 547 -29 581
rect -129 509 -29 547
rect 29 581 129 597
rect 29 547 45 581
rect 113 547 129 581
rect 29 509 129 547
rect 187 581 287 597
rect 187 547 203 581
rect 271 547 287 581
rect 187 509 287 547
rect 345 581 445 597
rect 345 547 361 581
rect 429 547 445 581
rect 345 509 445 547
rect 503 581 603 597
rect 503 547 519 581
rect 587 547 603 581
rect 503 509 603 547
rect 661 581 761 597
rect 661 547 677 581
rect 745 547 761 581
rect 661 509 761 547
rect 819 581 919 597
rect 819 547 835 581
rect 903 547 919 581
rect 819 509 919 547
rect 977 581 1077 597
rect 977 547 993 581
rect 1061 547 1077 581
rect 977 509 1077 547
rect 1135 581 1235 597
rect 1135 547 1151 581
rect 1219 547 1235 581
rect 1135 509 1235 547
rect -1235 71 -1135 109
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1235 21 -1135 37
rect -1077 71 -977 109
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 109
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 109
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 109
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 109
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 109
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 109
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 109
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 109
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 109
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect 1135 71 1235 109
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1135 21 1235 37
rect -1235 -37 -1135 -21
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1235 -109 -1135 -71
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -109 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -109 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -109 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -109 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -109 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -109 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -109 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -109 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -109 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -109 1077 -71
rect 1135 -37 1235 -21
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1135 -109 1235 -71
rect -1235 -547 -1135 -509
rect -1235 -581 -1219 -547
rect -1151 -581 -1135 -547
rect -1235 -597 -1135 -581
rect -1077 -547 -977 -509
rect -1077 -581 -1061 -547
rect -993 -581 -977 -547
rect -1077 -597 -977 -581
rect -919 -547 -819 -509
rect -919 -581 -903 -547
rect -835 -581 -819 -547
rect -919 -597 -819 -581
rect -761 -547 -661 -509
rect -761 -581 -745 -547
rect -677 -581 -661 -547
rect -761 -597 -661 -581
rect -603 -547 -503 -509
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -603 -597 -503 -581
rect -445 -547 -345 -509
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -445 -597 -345 -581
rect -287 -547 -187 -509
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -287 -597 -187 -581
rect -129 -547 -29 -509
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -509
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 29 -597 129 -581
rect 187 -547 287 -509
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 187 -597 287 -581
rect 345 -547 445 -509
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 345 -597 445 -581
rect 503 -547 603 -509
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 503 -597 603 -581
rect 661 -547 761 -509
rect 661 -581 677 -547
rect 745 -581 761 -547
rect 661 -597 761 -581
rect 819 -547 919 -509
rect 819 -581 835 -547
rect 903 -581 919 -547
rect 819 -597 919 -581
rect 977 -547 1077 -509
rect 977 -581 993 -547
rect 1061 -581 1077 -547
rect 977 -597 1077 -581
rect 1135 -547 1235 -509
rect 1135 -581 1151 -547
rect 1219 -581 1235 -547
rect 1135 -597 1235 -581
rect -1235 -655 -1135 -639
rect -1235 -689 -1219 -655
rect -1151 -689 -1135 -655
rect -1235 -727 -1135 -689
rect -1077 -655 -977 -639
rect -1077 -689 -1061 -655
rect -993 -689 -977 -655
rect -1077 -727 -977 -689
rect -919 -655 -819 -639
rect -919 -689 -903 -655
rect -835 -689 -819 -655
rect -919 -727 -819 -689
rect -761 -655 -661 -639
rect -761 -689 -745 -655
rect -677 -689 -661 -655
rect -761 -727 -661 -689
rect -603 -655 -503 -639
rect -603 -689 -587 -655
rect -519 -689 -503 -655
rect -603 -727 -503 -689
rect -445 -655 -345 -639
rect -445 -689 -429 -655
rect -361 -689 -345 -655
rect -445 -727 -345 -689
rect -287 -655 -187 -639
rect -287 -689 -271 -655
rect -203 -689 -187 -655
rect -287 -727 -187 -689
rect -129 -655 -29 -639
rect -129 -689 -113 -655
rect -45 -689 -29 -655
rect -129 -727 -29 -689
rect 29 -655 129 -639
rect 29 -689 45 -655
rect 113 -689 129 -655
rect 29 -727 129 -689
rect 187 -655 287 -639
rect 187 -689 203 -655
rect 271 -689 287 -655
rect 187 -727 287 -689
rect 345 -655 445 -639
rect 345 -689 361 -655
rect 429 -689 445 -655
rect 345 -727 445 -689
rect 503 -655 603 -639
rect 503 -689 519 -655
rect 587 -689 603 -655
rect 503 -727 603 -689
rect 661 -655 761 -639
rect 661 -689 677 -655
rect 745 -689 761 -655
rect 661 -727 761 -689
rect 819 -655 919 -639
rect 819 -689 835 -655
rect 903 -689 919 -655
rect 819 -727 919 -689
rect 977 -655 1077 -639
rect 977 -689 993 -655
rect 1061 -689 1077 -655
rect 977 -727 1077 -689
rect 1135 -655 1235 -639
rect 1135 -689 1151 -655
rect 1219 -689 1235 -655
rect 1135 -727 1235 -689
rect -1235 -1165 -1135 -1127
rect -1235 -1199 -1219 -1165
rect -1151 -1199 -1135 -1165
rect -1235 -1215 -1135 -1199
rect -1077 -1165 -977 -1127
rect -1077 -1199 -1061 -1165
rect -993 -1199 -977 -1165
rect -1077 -1215 -977 -1199
rect -919 -1165 -819 -1127
rect -919 -1199 -903 -1165
rect -835 -1199 -819 -1165
rect -919 -1215 -819 -1199
rect -761 -1165 -661 -1127
rect -761 -1199 -745 -1165
rect -677 -1199 -661 -1165
rect -761 -1215 -661 -1199
rect -603 -1165 -503 -1127
rect -603 -1199 -587 -1165
rect -519 -1199 -503 -1165
rect -603 -1215 -503 -1199
rect -445 -1165 -345 -1127
rect -445 -1199 -429 -1165
rect -361 -1199 -345 -1165
rect -445 -1215 -345 -1199
rect -287 -1165 -187 -1127
rect -287 -1199 -271 -1165
rect -203 -1199 -187 -1165
rect -287 -1215 -187 -1199
rect -129 -1165 -29 -1127
rect -129 -1199 -113 -1165
rect -45 -1199 -29 -1165
rect -129 -1215 -29 -1199
rect 29 -1165 129 -1127
rect 29 -1199 45 -1165
rect 113 -1199 129 -1165
rect 29 -1215 129 -1199
rect 187 -1165 287 -1127
rect 187 -1199 203 -1165
rect 271 -1199 287 -1165
rect 187 -1215 287 -1199
rect 345 -1165 445 -1127
rect 345 -1199 361 -1165
rect 429 -1199 445 -1165
rect 345 -1215 445 -1199
rect 503 -1165 603 -1127
rect 503 -1199 519 -1165
rect 587 -1199 603 -1165
rect 503 -1215 603 -1199
rect 661 -1165 761 -1127
rect 661 -1199 677 -1165
rect 745 -1199 761 -1165
rect 661 -1215 761 -1199
rect 819 -1165 919 -1127
rect 819 -1199 835 -1165
rect 903 -1199 919 -1165
rect 819 -1215 919 -1199
rect 977 -1165 1077 -1127
rect 977 -1199 993 -1165
rect 1061 -1199 1077 -1165
rect 977 -1215 1077 -1199
rect 1135 -1165 1235 -1127
rect 1135 -1199 1151 -1165
rect 1219 -1199 1235 -1165
rect 1135 -1215 1235 -1199
rect -1235 -1273 -1135 -1257
rect -1235 -1307 -1219 -1273
rect -1151 -1307 -1135 -1273
rect -1235 -1345 -1135 -1307
rect -1077 -1273 -977 -1257
rect -1077 -1307 -1061 -1273
rect -993 -1307 -977 -1273
rect -1077 -1345 -977 -1307
rect -919 -1273 -819 -1257
rect -919 -1307 -903 -1273
rect -835 -1307 -819 -1273
rect -919 -1345 -819 -1307
rect -761 -1273 -661 -1257
rect -761 -1307 -745 -1273
rect -677 -1307 -661 -1273
rect -761 -1345 -661 -1307
rect -603 -1273 -503 -1257
rect -603 -1307 -587 -1273
rect -519 -1307 -503 -1273
rect -603 -1345 -503 -1307
rect -445 -1273 -345 -1257
rect -445 -1307 -429 -1273
rect -361 -1307 -345 -1273
rect -445 -1345 -345 -1307
rect -287 -1273 -187 -1257
rect -287 -1307 -271 -1273
rect -203 -1307 -187 -1273
rect -287 -1345 -187 -1307
rect -129 -1273 -29 -1257
rect -129 -1307 -113 -1273
rect -45 -1307 -29 -1273
rect -129 -1345 -29 -1307
rect 29 -1273 129 -1257
rect 29 -1307 45 -1273
rect 113 -1307 129 -1273
rect 29 -1345 129 -1307
rect 187 -1273 287 -1257
rect 187 -1307 203 -1273
rect 271 -1307 287 -1273
rect 187 -1345 287 -1307
rect 345 -1273 445 -1257
rect 345 -1307 361 -1273
rect 429 -1307 445 -1273
rect 345 -1345 445 -1307
rect 503 -1273 603 -1257
rect 503 -1307 519 -1273
rect 587 -1307 603 -1273
rect 503 -1345 603 -1307
rect 661 -1273 761 -1257
rect 661 -1307 677 -1273
rect 745 -1307 761 -1273
rect 661 -1345 761 -1307
rect 819 -1273 919 -1257
rect 819 -1307 835 -1273
rect 903 -1307 919 -1273
rect 819 -1345 919 -1307
rect 977 -1273 1077 -1257
rect 977 -1307 993 -1273
rect 1061 -1307 1077 -1273
rect 977 -1345 1077 -1307
rect 1135 -1273 1235 -1257
rect 1135 -1307 1151 -1273
rect 1219 -1307 1235 -1273
rect 1135 -1345 1235 -1307
rect -1235 -1783 -1135 -1745
rect -1235 -1817 -1219 -1783
rect -1151 -1817 -1135 -1783
rect -1235 -1833 -1135 -1817
rect -1077 -1783 -977 -1745
rect -1077 -1817 -1061 -1783
rect -993 -1817 -977 -1783
rect -1077 -1833 -977 -1817
rect -919 -1783 -819 -1745
rect -919 -1817 -903 -1783
rect -835 -1817 -819 -1783
rect -919 -1833 -819 -1817
rect -761 -1783 -661 -1745
rect -761 -1817 -745 -1783
rect -677 -1817 -661 -1783
rect -761 -1833 -661 -1817
rect -603 -1783 -503 -1745
rect -603 -1817 -587 -1783
rect -519 -1817 -503 -1783
rect -603 -1833 -503 -1817
rect -445 -1783 -345 -1745
rect -445 -1817 -429 -1783
rect -361 -1817 -345 -1783
rect -445 -1833 -345 -1817
rect -287 -1783 -187 -1745
rect -287 -1817 -271 -1783
rect -203 -1817 -187 -1783
rect -287 -1833 -187 -1817
rect -129 -1783 -29 -1745
rect -129 -1817 -113 -1783
rect -45 -1817 -29 -1783
rect -129 -1833 -29 -1817
rect 29 -1783 129 -1745
rect 29 -1817 45 -1783
rect 113 -1817 129 -1783
rect 29 -1833 129 -1817
rect 187 -1783 287 -1745
rect 187 -1817 203 -1783
rect 271 -1817 287 -1783
rect 187 -1833 287 -1817
rect 345 -1783 445 -1745
rect 345 -1817 361 -1783
rect 429 -1817 445 -1783
rect 345 -1833 445 -1817
rect 503 -1783 603 -1745
rect 503 -1817 519 -1783
rect 587 -1817 603 -1783
rect 503 -1833 603 -1817
rect 661 -1783 761 -1745
rect 661 -1817 677 -1783
rect 745 -1817 761 -1783
rect 661 -1833 761 -1817
rect 819 -1783 919 -1745
rect 819 -1817 835 -1783
rect 903 -1817 919 -1783
rect 819 -1833 919 -1817
rect 977 -1783 1077 -1745
rect 977 -1817 993 -1783
rect 1061 -1817 1077 -1783
rect 977 -1833 1077 -1817
rect 1135 -1783 1235 -1745
rect 1135 -1817 1151 -1783
rect 1219 -1817 1235 -1783
rect 1135 -1833 1235 -1817
rect -1235 -1891 -1135 -1875
rect -1235 -1925 -1219 -1891
rect -1151 -1925 -1135 -1891
rect -1235 -1963 -1135 -1925
rect -1077 -1891 -977 -1875
rect -1077 -1925 -1061 -1891
rect -993 -1925 -977 -1891
rect -1077 -1963 -977 -1925
rect -919 -1891 -819 -1875
rect -919 -1925 -903 -1891
rect -835 -1925 -819 -1891
rect -919 -1963 -819 -1925
rect -761 -1891 -661 -1875
rect -761 -1925 -745 -1891
rect -677 -1925 -661 -1891
rect -761 -1963 -661 -1925
rect -603 -1891 -503 -1875
rect -603 -1925 -587 -1891
rect -519 -1925 -503 -1891
rect -603 -1963 -503 -1925
rect -445 -1891 -345 -1875
rect -445 -1925 -429 -1891
rect -361 -1925 -345 -1891
rect -445 -1963 -345 -1925
rect -287 -1891 -187 -1875
rect -287 -1925 -271 -1891
rect -203 -1925 -187 -1891
rect -287 -1963 -187 -1925
rect -129 -1891 -29 -1875
rect -129 -1925 -113 -1891
rect -45 -1925 -29 -1891
rect -129 -1963 -29 -1925
rect 29 -1891 129 -1875
rect 29 -1925 45 -1891
rect 113 -1925 129 -1891
rect 29 -1963 129 -1925
rect 187 -1891 287 -1875
rect 187 -1925 203 -1891
rect 271 -1925 287 -1891
rect 187 -1963 287 -1925
rect 345 -1891 445 -1875
rect 345 -1925 361 -1891
rect 429 -1925 445 -1891
rect 345 -1963 445 -1925
rect 503 -1891 603 -1875
rect 503 -1925 519 -1891
rect 587 -1925 603 -1891
rect 503 -1963 603 -1925
rect 661 -1891 761 -1875
rect 661 -1925 677 -1891
rect 745 -1925 761 -1891
rect 661 -1963 761 -1925
rect 819 -1891 919 -1875
rect 819 -1925 835 -1891
rect 903 -1925 919 -1891
rect 819 -1963 919 -1925
rect 977 -1891 1077 -1875
rect 977 -1925 993 -1891
rect 1061 -1925 1077 -1891
rect 977 -1963 1077 -1925
rect 1135 -1891 1235 -1875
rect 1135 -1925 1151 -1891
rect 1219 -1925 1235 -1891
rect 1135 -1963 1235 -1925
rect -1235 -2401 -1135 -2363
rect -1235 -2435 -1219 -2401
rect -1151 -2435 -1135 -2401
rect -1235 -2451 -1135 -2435
rect -1077 -2401 -977 -2363
rect -1077 -2435 -1061 -2401
rect -993 -2435 -977 -2401
rect -1077 -2451 -977 -2435
rect -919 -2401 -819 -2363
rect -919 -2435 -903 -2401
rect -835 -2435 -819 -2401
rect -919 -2451 -819 -2435
rect -761 -2401 -661 -2363
rect -761 -2435 -745 -2401
rect -677 -2435 -661 -2401
rect -761 -2451 -661 -2435
rect -603 -2401 -503 -2363
rect -603 -2435 -587 -2401
rect -519 -2435 -503 -2401
rect -603 -2451 -503 -2435
rect -445 -2401 -345 -2363
rect -445 -2435 -429 -2401
rect -361 -2435 -345 -2401
rect -445 -2451 -345 -2435
rect -287 -2401 -187 -2363
rect -287 -2435 -271 -2401
rect -203 -2435 -187 -2401
rect -287 -2451 -187 -2435
rect -129 -2401 -29 -2363
rect -129 -2435 -113 -2401
rect -45 -2435 -29 -2401
rect -129 -2451 -29 -2435
rect 29 -2401 129 -2363
rect 29 -2435 45 -2401
rect 113 -2435 129 -2401
rect 29 -2451 129 -2435
rect 187 -2401 287 -2363
rect 187 -2435 203 -2401
rect 271 -2435 287 -2401
rect 187 -2451 287 -2435
rect 345 -2401 445 -2363
rect 345 -2435 361 -2401
rect 429 -2435 445 -2401
rect 345 -2451 445 -2435
rect 503 -2401 603 -2363
rect 503 -2435 519 -2401
rect 587 -2435 603 -2401
rect 503 -2451 603 -2435
rect 661 -2401 761 -2363
rect 661 -2435 677 -2401
rect 745 -2435 761 -2401
rect 661 -2451 761 -2435
rect 819 -2401 919 -2363
rect 819 -2435 835 -2401
rect 903 -2435 919 -2401
rect 819 -2451 919 -2435
rect 977 -2401 1077 -2363
rect 977 -2435 993 -2401
rect 1061 -2435 1077 -2401
rect 977 -2451 1077 -2435
rect 1135 -2401 1235 -2363
rect 1135 -2435 1151 -2401
rect 1219 -2435 1235 -2401
rect 1135 -2451 1235 -2435
<< polycont >>
rect -1219 2401 -1151 2435
rect -1061 2401 -993 2435
rect -903 2401 -835 2435
rect -745 2401 -677 2435
rect -587 2401 -519 2435
rect -429 2401 -361 2435
rect -271 2401 -203 2435
rect -113 2401 -45 2435
rect 45 2401 113 2435
rect 203 2401 271 2435
rect 361 2401 429 2435
rect 519 2401 587 2435
rect 677 2401 745 2435
rect 835 2401 903 2435
rect 993 2401 1061 2435
rect 1151 2401 1219 2435
rect -1219 1891 -1151 1925
rect -1061 1891 -993 1925
rect -903 1891 -835 1925
rect -745 1891 -677 1925
rect -587 1891 -519 1925
rect -429 1891 -361 1925
rect -271 1891 -203 1925
rect -113 1891 -45 1925
rect 45 1891 113 1925
rect 203 1891 271 1925
rect 361 1891 429 1925
rect 519 1891 587 1925
rect 677 1891 745 1925
rect 835 1891 903 1925
rect 993 1891 1061 1925
rect 1151 1891 1219 1925
rect -1219 1783 -1151 1817
rect -1061 1783 -993 1817
rect -903 1783 -835 1817
rect -745 1783 -677 1817
rect -587 1783 -519 1817
rect -429 1783 -361 1817
rect -271 1783 -203 1817
rect -113 1783 -45 1817
rect 45 1783 113 1817
rect 203 1783 271 1817
rect 361 1783 429 1817
rect 519 1783 587 1817
rect 677 1783 745 1817
rect 835 1783 903 1817
rect 993 1783 1061 1817
rect 1151 1783 1219 1817
rect -1219 1273 -1151 1307
rect -1061 1273 -993 1307
rect -903 1273 -835 1307
rect -745 1273 -677 1307
rect -587 1273 -519 1307
rect -429 1273 -361 1307
rect -271 1273 -203 1307
rect -113 1273 -45 1307
rect 45 1273 113 1307
rect 203 1273 271 1307
rect 361 1273 429 1307
rect 519 1273 587 1307
rect 677 1273 745 1307
rect 835 1273 903 1307
rect 993 1273 1061 1307
rect 1151 1273 1219 1307
rect -1219 1165 -1151 1199
rect -1061 1165 -993 1199
rect -903 1165 -835 1199
rect -745 1165 -677 1199
rect -587 1165 -519 1199
rect -429 1165 -361 1199
rect -271 1165 -203 1199
rect -113 1165 -45 1199
rect 45 1165 113 1199
rect 203 1165 271 1199
rect 361 1165 429 1199
rect 519 1165 587 1199
rect 677 1165 745 1199
rect 835 1165 903 1199
rect 993 1165 1061 1199
rect 1151 1165 1219 1199
rect -1219 655 -1151 689
rect -1061 655 -993 689
rect -903 655 -835 689
rect -745 655 -677 689
rect -587 655 -519 689
rect -429 655 -361 689
rect -271 655 -203 689
rect -113 655 -45 689
rect 45 655 113 689
rect 203 655 271 689
rect 361 655 429 689
rect 519 655 587 689
rect 677 655 745 689
rect 835 655 903 689
rect 993 655 1061 689
rect 1151 655 1219 689
rect -1219 547 -1151 581
rect -1061 547 -993 581
rect -903 547 -835 581
rect -745 547 -677 581
rect -587 547 -519 581
rect -429 547 -361 581
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect 361 547 429 581
rect 519 547 587 581
rect 677 547 745 581
rect 835 547 903 581
rect 993 547 1061 581
rect 1151 547 1219 581
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect -1219 -581 -1151 -547
rect -1061 -581 -993 -547
rect -903 -581 -835 -547
rect -745 -581 -677 -547
rect -587 -581 -519 -547
rect -429 -581 -361 -547
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
rect 361 -581 429 -547
rect 519 -581 587 -547
rect 677 -581 745 -547
rect 835 -581 903 -547
rect 993 -581 1061 -547
rect 1151 -581 1219 -547
rect -1219 -689 -1151 -655
rect -1061 -689 -993 -655
rect -903 -689 -835 -655
rect -745 -689 -677 -655
rect -587 -689 -519 -655
rect -429 -689 -361 -655
rect -271 -689 -203 -655
rect -113 -689 -45 -655
rect 45 -689 113 -655
rect 203 -689 271 -655
rect 361 -689 429 -655
rect 519 -689 587 -655
rect 677 -689 745 -655
rect 835 -689 903 -655
rect 993 -689 1061 -655
rect 1151 -689 1219 -655
rect -1219 -1199 -1151 -1165
rect -1061 -1199 -993 -1165
rect -903 -1199 -835 -1165
rect -745 -1199 -677 -1165
rect -587 -1199 -519 -1165
rect -429 -1199 -361 -1165
rect -271 -1199 -203 -1165
rect -113 -1199 -45 -1165
rect 45 -1199 113 -1165
rect 203 -1199 271 -1165
rect 361 -1199 429 -1165
rect 519 -1199 587 -1165
rect 677 -1199 745 -1165
rect 835 -1199 903 -1165
rect 993 -1199 1061 -1165
rect 1151 -1199 1219 -1165
rect -1219 -1307 -1151 -1273
rect -1061 -1307 -993 -1273
rect -903 -1307 -835 -1273
rect -745 -1307 -677 -1273
rect -587 -1307 -519 -1273
rect -429 -1307 -361 -1273
rect -271 -1307 -203 -1273
rect -113 -1307 -45 -1273
rect 45 -1307 113 -1273
rect 203 -1307 271 -1273
rect 361 -1307 429 -1273
rect 519 -1307 587 -1273
rect 677 -1307 745 -1273
rect 835 -1307 903 -1273
rect 993 -1307 1061 -1273
rect 1151 -1307 1219 -1273
rect -1219 -1817 -1151 -1783
rect -1061 -1817 -993 -1783
rect -903 -1817 -835 -1783
rect -745 -1817 -677 -1783
rect -587 -1817 -519 -1783
rect -429 -1817 -361 -1783
rect -271 -1817 -203 -1783
rect -113 -1817 -45 -1783
rect 45 -1817 113 -1783
rect 203 -1817 271 -1783
rect 361 -1817 429 -1783
rect 519 -1817 587 -1783
rect 677 -1817 745 -1783
rect 835 -1817 903 -1783
rect 993 -1817 1061 -1783
rect 1151 -1817 1219 -1783
rect -1219 -1925 -1151 -1891
rect -1061 -1925 -993 -1891
rect -903 -1925 -835 -1891
rect -745 -1925 -677 -1891
rect -587 -1925 -519 -1891
rect -429 -1925 -361 -1891
rect -271 -1925 -203 -1891
rect -113 -1925 -45 -1891
rect 45 -1925 113 -1891
rect 203 -1925 271 -1891
rect 361 -1925 429 -1891
rect 519 -1925 587 -1891
rect 677 -1925 745 -1891
rect 835 -1925 903 -1891
rect 993 -1925 1061 -1891
rect 1151 -1925 1219 -1891
rect -1219 -2435 -1151 -2401
rect -1061 -2435 -993 -2401
rect -903 -2435 -835 -2401
rect -745 -2435 -677 -2401
rect -587 -2435 -519 -2401
rect -429 -2435 -361 -2401
rect -271 -2435 -203 -2401
rect -113 -2435 -45 -2401
rect 45 -2435 113 -2401
rect 203 -2435 271 -2401
rect 361 -2435 429 -2401
rect 519 -2435 587 -2401
rect 677 -2435 745 -2401
rect 835 -2435 903 -2401
rect 993 -2435 1061 -2401
rect 1151 -2435 1219 -2401
<< locali >>
rect -1395 2503 -1299 2537
rect 1299 2503 1395 2537
rect -1395 2441 -1361 2503
rect 1361 2441 1395 2503
rect -1235 2401 -1219 2435
rect -1151 2401 -1135 2435
rect -1077 2401 -1061 2435
rect -993 2401 -977 2435
rect -919 2401 -903 2435
rect -835 2401 -819 2435
rect -761 2401 -745 2435
rect -677 2401 -661 2435
rect -603 2401 -587 2435
rect -519 2401 -503 2435
rect -445 2401 -429 2435
rect -361 2401 -345 2435
rect -287 2401 -271 2435
rect -203 2401 -187 2435
rect -129 2401 -113 2435
rect -45 2401 -29 2435
rect 29 2401 45 2435
rect 113 2401 129 2435
rect 187 2401 203 2435
rect 271 2401 287 2435
rect 345 2401 361 2435
rect 429 2401 445 2435
rect 503 2401 519 2435
rect 587 2401 603 2435
rect 661 2401 677 2435
rect 745 2401 761 2435
rect 819 2401 835 2435
rect 903 2401 919 2435
rect 977 2401 993 2435
rect 1061 2401 1077 2435
rect 1135 2401 1151 2435
rect 1219 2401 1235 2435
rect -1281 2351 -1247 2367
rect -1281 1959 -1247 1975
rect -1123 2351 -1089 2367
rect -1123 1959 -1089 1975
rect -965 2351 -931 2367
rect -965 1959 -931 1975
rect -807 2351 -773 2367
rect -807 1959 -773 1975
rect -649 2351 -615 2367
rect -649 1959 -615 1975
rect -491 2351 -457 2367
rect -491 1959 -457 1975
rect -333 2351 -299 2367
rect -333 1959 -299 1975
rect -175 2351 -141 2367
rect -175 1959 -141 1975
rect -17 2351 17 2367
rect -17 1959 17 1975
rect 141 2351 175 2367
rect 141 1959 175 1975
rect 299 2351 333 2367
rect 299 1959 333 1975
rect 457 2351 491 2367
rect 457 1959 491 1975
rect 615 2351 649 2367
rect 615 1959 649 1975
rect 773 2351 807 2367
rect 773 1959 807 1975
rect 931 2351 965 2367
rect 931 1959 965 1975
rect 1089 2351 1123 2367
rect 1089 1959 1123 1975
rect 1247 2351 1281 2367
rect 1247 1959 1281 1975
rect -1235 1891 -1219 1925
rect -1151 1891 -1135 1925
rect -1077 1891 -1061 1925
rect -993 1891 -977 1925
rect -919 1891 -903 1925
rect -835 1891 -819 1925
rect -761 1891 -745 1925
rect -677 1891 -661 1925
rect -603 1891 -587 1925
rect -519 1891 -503 1925
rect -445 1891 -429 1925
rect -361 1891 -345 1925
rect -287 1891 -271 1925
rect -203 1891 -187 1925
rect -129 1891 -113 1925
rect -45 1891 -29 1925
rect 29 1891 45 1925
rect 113 1891 129 1925
rect 187 1891 203 1925
rect 271 1891 287 1925
rect 345 1891 361 1925
rect 429 1891 445 1925
rect 503 1891 519 1925
rect 587 1891 603 1925
rect 661 1891 677 1925
rect 745 1891 761 1925
rect 819 1891 835 1925
rect 903 1891 919 1925
rect 977 1891 993 1925
rect 1061 1891 1077 1925
rect 1135 1891 1151 1925
rect 1219 1891 1235 1925
rect -1235 1783 -1219 1817
rect -1151 1783 -1135 1817
rect -1077 1783 -1061 1817
rect -993 1783 -977 1817
rect -919 1783 -903 1817
rect -835 1783 -819 1817
rect -761 1783 -745 1817
rect -677 1783 -661 1817
rect -603 1783 -587 1817
rect -519 1783 -503 1817
rect -445 1783 -429 1817
rect -361 1783 -345 1817
rect -287 1783 -271 1817
rect -203 1783 -187 1817
rect -129 1783 -113 1817
rect -45 1783 -29 1817
rect 29 1783 45 1817
rect 113 1783 129 1817
rect 187 1783 203 1817
rect 271 1783 287 1817
rect 345 1783 361 1817
rect 429 1783 445 1817
rect 503 1783 519 1817
rect 587 1783 603 1817
rect 661 1783 677 1817
rect 745 1783 761 1817
rect 819 1783 835 1817
rect 903 1783 919 1817
rect 977 1783 993 1817
rect 1061 1783 1077 1817
rect 1135 1783 1151 1817
rect 1219 1783 1235 1817
rect -1281 1733 -1247 1749
rect -1281 1341 -1247 1357
rect -1123 1733 -1089 1749
rect -1123 1341 -1089 1357
rect -965 1733 -931 1749
rect -965 1341 -931 1357
rect -807 1733 -773 1749
rect -807 1341 -773 1357
rect -649 1733 -615 1749
rect -649 1341 -615 1357
rect -491 1733 -457 1749
rect -491 1341 -457 1357
rect -333 1733 -299 1749
rect -333 1341 -299 1357
rect -175 1733 -141 1749
rect -175 1341 -141 1357
rect -17 1733 17 1749
rect -17 1341 17 1357
rect 141 1733 175 1749
rect 141 1341 175 1357
rect 299 1733 333 1749
rect 299 1341 333 1357
rect 457 1733 491 1749
rect 457 1341 491 1357
rect 615 1733 649 1749
rect 615 1341 649 1357
rect 773 1733 807 1749
rect 773 1341 807 1357
rect 931 1733 965 1749
rect 931 1341 965 1357
rect 1089 1733 1123 1749
rect 1089 1341 1123 1357
rect 1247 1733 1281 1749
rect 1247 1341 1281 1357
rect -1235 1273 -1219 1307
rect -1151 1273 -1135 1307
rect -1077 1273 -1061 1307
rect -993 1273 -977 1307
rect -919 1273 -903 1307
rect -835 1273 -819 1307
rect -761 1273 -745 1307
rect -677 1273 -661 1307
rect -603 1273 -587 1307
rect -519 1273 -503 1307
rect -445 1273 -429 1307
rect -361 1273 -345 1307
rect -287 1273 -271 1307
rect -203 1273 -187 1307
rect -129 1273 -113 1307
rect -45 1273 -29 1307
rect 29 1273 45 1307
rect 113 1273 129 1307
rect 187 1273 203 1307
rect 271 1273 287 1307
rect 345 1273 361 1307
rect 429 1273 445 1307
rect 503 1273 519 1307
rect 587 1273 603 1307
rect 661 1273 677 1307
rect 745 1273 761 1307
rect 819 1273 835 1307
rect 903 1273 919 1307
rect 977 1273 993 1307
rect 1061 1273 1077 1307
rect 1135 1273 1151 1307
rect 1219 1273 1235 1307
rect -1235 1165 -1219 1199
rect -1151 1165 -1135 1199
rect -1077 1165 -1061 1199
rect -993 1165 -977 1199
rect -919 1165 -903 1199
rect -835 1165 -819 1199
rect -761 1165 -745 1199
rect -677 1165 -661 1199
rect -603 1165 -587 1199
rect -519 1165 -503 1199
rect -445 1165 -429 1199
rect -361 1165 -345 1199
rect -287 1165 -271 1199
rect -203 1165 -187 1199
rect -129 1165 -113 1199
rect -45 1165 -29 1199
rect 29 1165 45 1199
rect 113 1165 129 1199
rect 187 1165 203 1199
rect 271 1165 287 1199
rect 345 1165 361 1199
rect 429 1165 445 1199
rect 503 1165 519 1199
rect 587 1165 603 1199
rect 661 1165 677 1199
rect 745 1165 761 1199
rect 819 1165 835 1199
rect 903 1165 919 1199
rect 977 1165 993 1199
rect 1061 1165 1077 1199
rect 1135 1165 1151 1199
rect 1219 1165 1235 1199
rect -1281 1115 -1247 1131
rect -1281 723 -1247 739
rect -1123 1115 -1089 1131
rect -1123 723 -1089 739
rect -965 1115 -931 1131
rect -965 723 -931 739
rect -807 1115 -773 1131
rect -807 723 -773 739
rect -649 1115 -615 1131
rect -649 723 -615 739
rect -491 1115 -457 1131
rect -491 723 -457 739
rect -333 1115 -299 1131
rect -333 723 -299 739
rect -175 1115 -141 1131
rect -175 723 -141 739
rect -17 1115 17 1131
rect -17 723 17 739
rect 141 1115 175 1131
rect 141 723 175 739
rect 299 1115 333 1131
rect 299 723 333 739
rect 457 1115 491 1131
rect 457 723 491 739
rect 615 1115 649 1131
rect 615 723 649 739
rect 773 1115 807 1131
rect 773 723 807 739
rect 931 1115 965 1131
rect 931 723 965 739
rect 1089 1115 1123 1131
rect 1089 723 1123 739
rect 1247 1115 1281 1131
rect 1247 723 1281 739
rect -1235 655 -1219 689
rect -1151 655 -1135 689
rect -1077 655 -1061 689
rect -993 655 -977 689
rect -919 655 -903 689
rect -835 655 -819 689
rect -761 655 -745 689
rect -677 655 -661 689
rect -603 655 -587 689
rect -519 655 -503 689
rect -445 655 -429 689
rect -361 655 -345 689
rect -287 655 -271 689
rect -203 655 -187 689
rect -129 655 -113 689
rect -45 655 -29 689
rect 29 655 45 689
rect 113 655 129 689
rect 187 655 203 689
rect 271 655 287 689
rect 345 655 361 689
rect 429 655 445 689
rect 503 655 519 689
rect 587 655 603 689
rect 661 655 677 689
rect 745 655 761 689
rect 819 655 835 689
rect 903 655 919 689
rect 977 655 993 689
rect 1061 655 1077 689
rect 1135 655 1151 689
rect 1219 655 1235 689
rect -1235 547 -1219 581
rect -1151 547 -1135 581
rect -1077 547 -1061 581
rect -993 547 -977 581
rect -919 547 -903 581
rect -835 547 -819 581
rect -761 547 -745 581
rect -677 547 -661 581
rect -603 547 -587 581
rect -519 547 -503 581
rect -445 547 -429 581
rect -361 547 -345 581
rect -287 547 -271 581
rect -203 547 -187 581
rect -129 547 -113 581
rect -45 547 -29 581
rect 29 547 45 581
rect 113 547 129 581
rect 187 547 203 581
rect 271 547 287 581
rect 345 547 361 581
rect 429 547 445 581
rect 503 547 519 581
rect 587 547 603 581
rect 661 547 677 581
rect 745 547 761 581
rect 819 547 835 581
rect 903 547 919 581
rect 977 547 993 581
rect 1061 547 1077 581
rect 1135 547 1151 581
rect 1219 547 1235 581
rect -1281 497 -1247 513
rect -1281 105 -1247 121
rect -1123 497 -1089 513
rect -1123 105 -1089 121
rect -965 497 -931 513
rect -965 105 -931 121
rect -807 497 -773 513
rect -807 105 -773 121
rect -649 497 -615 513
rect -649 105 -615 121
rect -491 497 -457 513
rect -491 105 -457 121
rect -333 497 -299 513
rect -333 105 -299 121
rect -175 497 -141 513
rect -175 105 -141 121
rect -17 497 17 513
rect -17 105 17 121
rect 141 497 175 513
rect 141 105 175 121
rect 299 497 333 513
rect 299 105 333 121
rect 457 497 491 513
rect 457 105 491 121
rect 615 497 649 513
rect 615 105 649 121
rect 773 497 807 513
rect 773 105 807 121
rect 931 497 965 513
rect 931 105 965 121
rect 1089 497 1123 513
rect 1089 105 1123 121
rect 1247 497 1281 513
rect 1247 105 1281 121
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect 1135 37 1151 71
rect 1219 37 1235 71
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect -1281 -121 -1247 -105
rect -1281 -513 -1247 -497
rect -1123 -121 -1089 -105
rect -1123 -513 -1089 -497
rect -965 -121 -931 -105
rect -965 -513 -931 -497
rect -807 -121 -773 -105
rect -807 -513 -773 -497
rect -649 -121 -615 -105
rect -649 -513 -615 -497
rect -491 -121 -457 -105
rect -491 -513 -457 -497
rect -333 -121 -299 -105
rect -333 -513 -299 -497
rect -175 -121 -141 -105
rect -175 -513 -141 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 141 -121 175 -105
rect 141 -513 175 -497
rect 299 -121 333 -105
rect 299 -513 333 -497
rect 457 -121 491 -105
rect 457 -513 491 -497
rect 615 -121 649 -105
rect 615 -513 649 -497
rect 773 -121 807 -105
rect 773 -513 807 -497
rect 931 -121 965 -105
rect 931 -513 965 -497
rect 1089 -121 1123 -105
rect 1089 -513 1123 -497
rect 1247 -121 1281 -105
rect 1247 -513 1281 -497
rect -1235 -581 -1219 -547
rect -1151 -581 -1135 -547
rect -1077 -581 -1061 -547
rect -993 -581 -977 -547
rect -919 -581 -903 -547
rect -835 -581 -819 -547
rect -761 -581 -745 -547
rect -677 -581 -661 -547
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 661 -581 677 -547
rect 745 -581 761 -547
rect 819 -581 835 -547
rect 903 -581 919 -547
rect 977 -581 993 -547
rect 1061 -581 1077 -547
rect 1135 -581 1151 -547
rect 1219 -581 1235 -547
rect -1235 -689 -1219 -655
rect -1151 -689 -1135 -655
rect -1077 -689 -1061 -655
rect -993 -689 -977 -655
rect -919 -689 -903 -655
rect -835 -689 -819 -655
rect -761 -689 -745 -655
rect -677 -689 -661 -655
rect -603 -689 -587 -655
rect -519 -689 -503 -655
rect -445 -689 -429 -655
rect -361 -689 -345 -655
rect -287 -689 -271 -655
rect -203 -689 -187 -655
rect -129 -689 -113 -655
rect -45 -689 -29 -655
rect 29 -689 45 -655
rect 113 -689 129 -655
rect 187 -689 203 -655
rect 271 -689 287 -655
rect 345 -689 361 -655
rect 429 -689 445 -655
rect 503 -689 519 -655
rect 587 -689 603 -655
rect 661 -689 677 -655
rect 745 -689 761 -655
rect 819 -689 835 -655
rect 903 -689 919 -655
rect 977 -689 993 -655
rect 1061 -689 1077 -655
rect 1135 -689 1151 -655
rect 1219 -689 1235 -655
rect -1281 -739 -1247 -723
rect -1281 -1131 -1247 -1115
rect -1123 -739 -1089 -723
rect -1123 -1131 -1089 -1115
rect -965 -739 -931 -723
rect -965 -1131 -931 -1115
rect -807 -739 -773 -723
rect -807 -1131 -773 -1115
rect -649 -739 -615 -723
rect -649 -1131 -615 -1115
rect -491 -739 -457 -723
rect -491 -1131 -457 -1115
rect -333 -739 -299 -723
rect -333 -1131 -299 -1115
rect -175 -739 -141 -723
rect -175 -1131 -141 -1115
rect -17 -739 17 -723
rect -17 -1131 17 -1115
rect 141 -739 175 -723
rect 141 -1131 175 -1115
rect 299 -739 333 -723
rect 299 -1131 333 -1115
rect 457 -739 491 -723
rect 457 -1131 491 -1115
rect 615 -739 649 -723
rect 615 -1131 649 -1115
rect 773 -739 807 -723
rect 773 -1131 807 -1115
rect 931 -739 965 -723
rect 931 -1131 965 -1115
rect 1089 -739 1123 -723
rect 1089 -1131 1123 -1115
rect 1247 -739 1281 -723
rect 1247 -1131 1281 -1115
rect -1235 -1199 -1219 -1165
rect -1151 -1199 -1135 -1165
rect -1077 -1199 -1061 -1165
rect -993 -1199 -977 -1165
rect -919 -1199 -903 -1165
rect -835 -1199 -819 -1165
rect -761 -1199 -745 -1165
rect -677 -1199 -661 -1165
rect -603 -1199 -587 -1165
rect -519 -1199 -503 -1165
rect -445 -1199 -429 -1165
rect -361 -1199 -345 -1165
rect -287 -1199 -271 -1165
rect -203 -1199 -187 -1165
rect -129 -1199 -113 -1165
rect -45 -1199 -29 -1165
rect 29 -1199 45 -1165
rect 113 -1199 129 -1165
rect 187 -1199 203 -1165
rect 271 -1199 287 -1165
rect 345 -1199 361 -1165
rect 429 -1199 445 -1165
rect 503 -1199 519 -1165
rect 587 -1199 603 -1165
rect 661 -1199 677 -1165
rect 745 -1199 761 -1165
rect 819 -1199 835 -1165
rect 903 -1199 919 -1165
rect 977 -1199 993 -1165
rect 1061 -1199 1077 -1165
rect 1135 -1199 1151 -1165
rect 1219 -1199 1235 -1165
rect -1235 -1307 -1219 -1273
rect -1151 -1307 -1135 -1273
rect -1077 -1307 -1061 -1273
rect -993 -1307 -977 -1273
rect -919 -1307 -903 -1273
rect -835 -1307 -819 -1273
rect -761 -1307 -745 -1273
rect -677 -1307 -661 -1273
rect -603 -1307 -587 -1273
rect -519 -1307 -503 -1273
rect -445 -1307 -429 -1273
rect -361 -1307 -345 -1273
rect -287 -1307 -271 -1273
rect -203 -1307 -187 -1273
rect -129 -1307 -113 -1273
rect -45 -1307 -29 -1273
rect 29 -1307 45 -1273
rect 113 -1307 129 -1273
rect 187 -1307 203 -1273
rect 271 -1307 287 -1273
rect 345 -1307 361 -1273
rect 429 -1307 445 -1273
rect 503 -1307 519 -1273
rect 587 -1307 603 -1273
rect 661 -1307 677 -1273
rect 745 -1307 761 -1273
rect 819 -1307 835 -1273
rect 903 -1307 919 -1273
rect 977 -1307 993 -1273
rect 1061 -1307 1077 -1273
rect 1135 -1307 1151 -1273
rect 1219 -1307 1235 -1273
rect -1281 -1357 -1247 -1341
rect -1281 -1749 -1247 -1733
rect -1123 -1357 -1089 -1341
rect -1123 -1749 -1089 -1733
rect -965 -1357 -931 -1341
rect -965 -1749 -931 -1733
rect -807 -1357 -773 -1341
rect -807 -1749 -773 -1733
rect -649 -1357 -615 -1341
rect -649 -1749 -615 -1733
rect -491 -1357 -457 -1341
rect -491 -1749 -457 -1733
rect -333 -1357 -299 -1341
rect -333 -1749 -299 -1733
rect -175 -1357 -141 -1341
rect -175 -1749 -141 -1733
rect -17 -1357 17 -1341
rect -17 -1749 17 -1733
rect 141 -1357 175 -1341
rect 141 -1749 175 -1733
rect 299 -1357 333 -1341
rect 299 -1749 333 -1733
rect 457 -1357 491 -1341
rect 457 -1749 491 -1733
rect 615 -1357 649 -1341
rect 615 -1749 649 -1733
rect 773 -1357 807 -1341
rect 773 -1749 807 -1733
rect 931 -1357 965 -1341
rect 931 -1749 965 -1733
rect 1089 -1357 1123 -1341
rect 1089 -1749 1123 -1733
rect 1247 -1357 1281 -1341
rect 1247 -1749 1281 -1733
rect -1235 -1817 -1219 -1783
rect -1151 -1817 -1135 -1783
rect -1077 -1817 -1061 -1783
rect -993 -1817 -977 -1783
rect -919 -1817 -903 -1783
rect -835 -1817 -819 -1783
rect -761 -1817 -745 -1783
rect -677 -1817 -661 -1783
rect -603 -1817 -587 -1783
rect -519 -1817 -503 -1783
rect -445 -1817 -429 -1783
rect -361 -1817 -345 -1783
rect -287 -1817 -271 -1783
rect -203 -1817 -187 -1783
rect -129 -1817 -113 -1783
rect -45 -1817 -29 -1783
rect 29 -1817 45 -1783
rect 113 -1817 129 -1783
rect 187 -1817 203 -1783
rect 271 -1817 287 -1783
rect 345 -1817 361 -1783
rect 429 -1817 445 -1783
rect 503 -1817 519 -1783
rect 587 -1817 603 -1783
rect 661 -1817 677 -1783
rect 745 -1817 761 -1783
rect 819 -1817 835 -1783
rect 903 -1817 919 -1783
rect 977 -1817 993 -1783
rect 1061 -1817 1077 -1783
rect 1135 -1817 1151 -1783
rect 1219 -1817 1235 -1783
rect -1235 -1925 -1219 -1891
rect -1151 -1925 -1135 -1891
rect -1077 -1925 -1061 -1891
rect -993 -1925 -977 -1891
rect -919 -1925 -903 -1891
rect -835 -1925 -819 -1891
rect -761 -1925 -745 -1891
rect -677 -1925 -661 -1891
rect -603 -1925 -587 -1891
rect -519 -1925 -503 -1891
rect -445 -1925 -429 -1891
rect -361 -1925 -345 -1891
rect -287 -1925 -271 -1891
rect -203 -1925 -187 -1891
rect -129 -1925 -113 -1891
rect -45 -1925 -29 -1891
rect 29 -1925 45 -1891
rect 113 -1925 129 -1891
rect 187 -1925 203 -1891
rect 271 -1925 287 -1891
rect 345 -1925 361 -1891
rect 429 -1925 445 -1891
rect 503 -1925 519 -1891
rect 587 -1925 603 -1891
rect 661 -1925 677 -1891
rect 745 -1925 761 -1891
rect 819 -1925 835 -1891
rect 903 -1925 919 -1891
rect 977 -1925 993 -1891
rect 1061 -1925 1077 -1891
rect 1135 -1925 1151 -1891
rect 1219 -1925 1235 -1891
rect -1281 -1975 -1247 -1959
rect -1281 -2367 -1247 -2351
rect -1123 -1975 -1089 -1959
rect -1123 -2367 -1089 -2351
rect -965 -1975 -931 -1959
rect -965 -2367 -931 -2351
rect -807 -1975 -773 -1959
rect -807 -2367 -773 -2351
rect -649 -1975 -615 -1959
rect -649 -2367 -615 -2351
rect -491 -1975 -457 -1959
rect -491 -2367 -457 -2351
rect -333 -1975 -299 -1959
rect -333 -2367 -299 -2351
rect -175 -1975 -141 -1959
rect -175 -2367 -141 -2351
rect -17 -1975 17 -1959
rect -17 -2367 17 -2351
rect 141 -1975 175 -1959
rect 141 -2367 175 -2351
rect 299 -1975 333 -1959
rect 299 -2367 333 -2351
rect 457 -1975 491 -1959
rect 457 -2367 491 -2351
rect 615 -1975 649 -1959
rect 615 -2367 649 -2351
rect 773 -1975 807 -1959
rect 773 -2367 807 -2351
rect 931 -1975 965 -1959
rect 931 -2367 965 -2351
rect 1089 -1975 1123 -1959
rect 1089 -2367 1123 -2351
rect 1247 -1975 1281 -1959
rect 1247 -2367 1281 -2351
rect -1235 -2435 -1219 -2401
rect -1151 -2435 -1135 -2401
rect -1077 -2435 -1061 -2401
rect -993 -2435 -977 -2401
rect -919 -2435 -903 -2401
rect -835 -2435 -819 -2401
rect -761 -2435 -745 -2401
rect -677 -2435 -661 -2401
rect -603 -2435 -587 -2401
rect -519 -2435 -503 -2401
rect -445 -2435 -429 -2401
rect -361 -2435 -345 -2401
rect -287 -2435 -271 -2401
rect -203 -2435 -187 -2401
rect -129 -2435 -113 -2401
rect -45 -2435 -29 -2401
rect 29 -2435 45 -2401
rect 113 -2435 129 -2401
rect 187 -2435 203 -2401
rect 271 -2435 287 -2401
rect 345 -2435 361 -2401
rect 429 -2435 445 -2401
rect 503 -2435 519 -2401
rect 587 -2435 603 -2401
rect 661 -2435 677 -2401
rect 745 -2435 761 -2401
rect 819 -2435 835 -2401
rect 903 -2435 919 -2401
rect 977 -2435 993 -2401
rect 1061 -2435 1077 -2401
rect 1135 -2435 1151 -2401
rect 1219 -2435 1235 -2401
rect -1395 -2503 -1361 -2441
rect 1361 -2503 1395 -2441
rect -1395 -2537 -1299 -2503
rect 1299 -2537 1395 -2503
<< viali >>
rect -1219 2401 -1151 2435
rect -1061 2401 -993 2435
rect -903 2401 -835 2435
rect -745 2401 -677 2435
rect -587 2401 -519 2435
rect -429 2401 -361 2435
rect -271 2401 -203 2435
rect -113 2401 -45 2435
rect 45 2401 113 2435
rect 203 2401 271 2435
rect 361 2401 429 2435
rect 519 2401 587 2435
rect 677 2401 745 2435
rect 835 2401 903 2435
rect 993 2401 1061 2435
rect 1151 2401 1219 2435
rect -1281 1975 -1247 2351
rect -1123 1975 -1089 2351
rect -965 1975 -931 2351
rect -807 1975 -773 2351
rect -649 1975 -615 2351
rect -491 1975 -457 2351
rect -333 1975 -299 2351
rect -175 1975 -141 2351
rect -17 1975 17 2351
rect 141 1975 175 2351
rect 299 1975 333 2351
rect 457 1975 491 2351
rect 615 1975 649 2351
rect 773 1975 807 2351
rect 931 1975 965 2351
rect 1089 1975 1123 2351
rect 1247 1975 1281 2351
rect -1219 1891 -1151 1925
rect -1061 1891 -993 1925
rect -903 1891 -835 1925
rect -745 1891 -677 1925
rect -587 1891 -519 1925
rect -429 1891 -361 1925
rect -271 1891 -203 1925
rect -113 1891 -45 1925
rect 45 1891 113 1925
rect 203 1891 271 1925
rect 361 1891 429 1925
rect 519 1891 587 1925
rect 677 1891 745 1925
rect 835 1891 903 1925
rect 993 1891 1061 1925
rect 1151 1891 1219 1925
rect -1219 1783 -1151 1817
rect -1061 1783 -993 1817
rect -903 1783 -835 1817
rect -745 1783 -677 1817
rect -587 1783 -519 1817
rect -429 1783 -361 1817
rect -271 1783 -203 1817
rect -113 1783 -45 1817
rect 45 1783 113 1817
rect 203 1783 271 1817
rect 361 1783 429 1817
rect 519 1783 587 1817
rect 677 1783 745 1817
rect 835 1783 903 1817
rect 993 1783 1061 1817
rect 1151 1783 1219 1817
rect -1281 1357 -1247 1733
rect -1123 1357 -1089 1733
rect -965 1357 -931 1733
rect -807 1357 -773 1733
rect -649 1357 -615 1733
rect -491 1357 -457 1733
rect -333 1357 -299 1733
rect -175 1357 -141 1733
rect -17 1357 17 1733
rect 141 1357 175 1733
rect 299 1357 333 1733
rect 457 1357 491 1733
rect 615 1357 649 1733
rect 773 1357 807 1733
rect 931 1357 965 1733
rect 1089 1357 1123 1733
rect 1247 1357 1281 1733
rect -1219 1273 -1151 1307
rect -1061 1273 -993 1307
rect -903 1273 -835 1307
rect -745 1273 -677 1307
rect -587 1273 -519 1307
rect -429 1273 -361 1307
rect -271 1273 -203 1307
rect -113 1273 -45 1307
rect 45 1273 113 1307
rect 203 1273 271 1307
rect 361 1273 429 1307
rect 519 1273 587 1307
rect 677 1273 745 1307
rect 835 1273 903 1307
rect 993 1273 1061 1307
rect 1151 1273 1219 1307
rect -1219 1165 -1151 1199
rect -1061 1165 -993 1199
rect -903 1165 -835 1199
rect -745 1165 -677 1199
rect -587 1165 -519 1199
rect -429 1165 -361 1199
rect -271 1165 -203 1199
rect -113 1165 -45 1199
rect 45 1165 113 1199
rect 203 1165 271 1199
rect 361 1165 429 1199
rect 519 1165 587 1199
rect 677 1165 745 1199
rect 835 1165 903 1199
rect 993 1165 1061 1199
rect 1151 1165 1219 1199
rect -1281 739 -1247 1115
rect -1123 739 -1089 1115
rect -965 739 -931 1115
rect -807 739 -773 1115
rect -649 739 -615 1115
rect -491 739 -457 1115
rect -333 739 -299 1115
rect -175 739 -141 1115
rect -17 739 17 1115
rect 141 739 175 1115
rect 299 739 333 1115
rect 457 739 491 1115
rect 615 739 649 1115
rect 773 739 807 1115
rect 931 739 965 1115
rect 1089 739 1123 1115
rect 1247 739 1281 1115
rect -1219 655 -1151 689
rect -1061 655 -993 689
rect -903 655 -835 689
rect -745 655 -677 689
rect -587 655 -519 689
rect -429 655 -361 689
rect -271 655 -203 689
rect -113 655 -45 689
rect 45 655 113 689
rect 203 655 271 689
rect 361 655 429 689
rect 519 655 587 689
rect 677 655 745 689
rect 835 655 903 689
rect 993 655 1061 689
rect 1151 655 1219 689
rect -1219 547 -1151 581
rect -1061 547 -993 581
rect -903 547 -835 581
rect -745 547 -677 581
rect -587 547 -519 581
rect -429 547 -361 581
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect 361 547 429 581
rect 519 547 587 581
rect 677 547 745 581
rect 835 547 903 581
rect 993 547 1061 581
rect 1151 547 1219 581
rect -1281 121 -1247 497
rect -1123 121 -1089 497
rect -965 121 -931 497
rect -807 121 -773 497
rect -649 121 -615 497
rect -491 121 -457 497
rect -333 121 -299 497
rect -175 121 -141 497
rect -17 121 17 497
rect 141 121 175 497
rect 299 121 333 497
rect 457 121 491 497
rect 615 121 649 497
rect 773 121 807 497
rect 931 121 965 497
rect 1089 121 1123 497
rect 1247 121 1281 497
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect -1281 -497 -1247 -121
rect -1123 -497 -1089 -121
rect -965 -497 -931 -121
rect -807 -497 -773 -121
rect -649 -497 -615 -121
rect -491 -497 -457 -121
rect -333 -497 -299 -121
rect -175 -497 -141 -121
rect -17 -497 17 -121
rect 141 -497 175 -121
rect 299 -497 333 -121
rect 457 -497 491 -121
rect 615 -497 649 -121
rect 773 -497 807 -121
rect 931 -497 965 -121
rect 1089 -497 1123 -121
rect 1247 -497 1281 -121
rect -1219 -581 -1151 -547
rect -1061 -581 -993 -547
rect -903 -581 -835 -547
rect -745 -581 -677 -547
rect -587 -581 -519 -547
rect -429 -581 -361 -547
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
rect 361 -581 429 -547
rect 519 -581 587 -547
rect 677 -581 745 -547
rect 835 -581 903 -547
rect 993 -581 1061 -547
rect 1151 -581 1219 -547
rect -1219 -689 -1151 -655
rect -1061 -689 -993 -655
rect -903 -689 -835 -655
rect -745 -689 -677 -655
rect -587 -689 -519 -655
rect -429 -689 -361 -655
rect -271 -689 -203 -655
rect -113 -689 -45 -655
rect 45 -689 113 -655
rect 203 -689 271 -655
rect 361 -689 429 -655
rect 519 -689 587 -655
rect 677 -689 745 -655
rect 835 -689 903 -655
rect 993 -689 1061 -655
rect 1151 -689 1219 -655
rect -1281 -1115 -1247 -739
rect -1123 -1115 -1089 -739
rect -965 -1115 -931 -739
rect -807 -1115 -773 -739
rect -649 -1115 -615 -739
rect -491 -1115 -457 -739
rect -333 -1115 -299 -739
rect -175 -1115 -141 -739
rect -17 -1115 17 -739
rect 141 -1115 175 -739
rect 299 -1115 333 -739
rect 457 -1115 491 -739
rect 615 -1115 649 -739
rect 773 -1115 807 -739
rect 931 -1115 965 -739
rect 1089 -1115 1123 -739
rect 1247 -1115 1281 -739
rect -1219 -1199 -1151 -1165
rect -1061 -1199 -993 -1165
rect -903 -1199 -835 -1165
rect -745 -1199 -677 -1165
rect -587 -1199 -519 -1165
rect -429 -1199 -361 -1165
rect -271 -1199 -203 -1165
rect -113 -1199 -45 -1165
rect 45 -1199 113 -1165
rect 203 -1199 271 -1165
rect 361 -1199 429 -1165
rect 519 -1199 587 -1165
rect 677 -1199 745 -1165
rect 835 -1199 903 -1165
rect 993 -1199 1061 -1165
rect 1151 -1199 1219 -1165
rect -1219 -1307 -1151 -1273
rect -1061 -1307 -993 -1273
rect -903 -1307 -835 -1273
rect -745 -1307 -677 -1273
rect -587 -1307 -519 -1273
rect -429 -1307 -361 -1273
rect -271 -1307 -203 -1273
rect -113 -1307 -45 -1273
rect 45 -1307 113 -1273
rect 203 -1307 271 -1273
rect 361 -1307 429 -1273
rect 519 -1307 587 -1273
rect 677 -1307 745 -1273
rect 835 -1307 903 -1273
rect 993 -1307 1061 -1273
rect 1151 -1307 1219 -1273
rect -1281 -1733 -1247 -1357
rect -1123 -1733 -1089 -1357
rect -965 -1733 -931 -1357
rect -807 -1733 -773 -1357
rect -649 -1733 -615 -1357
rect -491 -1733 -457 -1357
rect -333 -1733 -299 -1357
rect -175 -1733 -141 -1357
rect -17 -1733 17 -1357
rect 141 -1733 175 -1357
rect 299 -1733 333 -1357
rect 457 -1733 491 -1357
rect 615 -1733 649 -1357
rect 773 -1733 807 -1357
rect 931 -1733 965 -1357
rect 1089 -1733 1123 -1357
rect 1247 -1733 1281 -1357
rect -1219 -1817 -1151 -1783
rect -1061 -1817 -993 -1783
rect -903 -1817 -835 -1783
rect -745 -1817 -677 -1783
rect -587 -1817 -519 -1783
rect -429 -1817 -361 -1783
rect -271 -1817 -203 -1783
rect -113 -1817 -45 -1783
rect 45 -1817 113 -1783
rect 203 -1817 271 -1783
rect 361 -1817 429 -1783
rect 519 -1817 587 -1783
rect 677 -1817 745 -1783
rect 835 -1817 903 -1783
rect 993 -1817 1061 -1783
rect 1151 -1817 1219 -1783
rect -1219 -1925 -1151 -1891
rect -1061 -1925 -993 -1891
rect -903 -1925 -835 -1891
rect -745 -1925 -677 -1891
rect -587 -1925 -519 -1891
rect -429 -1925 -361 -1891
rect -271 -1925 -203 -1891
rect -113 -1925 -45 -1891
rect 45 -1925 113 -1891
rect 203 -1925 271 -1891
rect 361 -1925 429 -1891
rect 519 -1925 587 -1891
rect 677 -1925 745 -1891
rect 835 -1925 903 -1891
rect 993 -1925 1061 -1891
rect 1151 -1925 1219 -1891
rect -1281 -2351 -1247 -1975
rect -1123 -2351 -1089 -1975
rect -965 -2351 -931 -1975
rect -807 -2351 -773 -1975
rect -649 -2351 -615 -1975
rect -491 -2351 -457 -1975
rect -333 -2351 -299 -1975
rect -175 -2351 -141 -1975
rect -17 -2351 17 -1975
rect 141 -2351 175 -1975
rect 299 -2351 333 -1975
rect 457 -2351 491 -1975
rect 615 -2351 649 -1975
rect 773 -2351 807 -1975
rect 931 -2351 965 -1975
rect 1089 -2351 1123 -1975
rect 1247 -2351 1281 -1975
rect -1219 -2435 -1151 -2401
rect -1061 -2435 -993 -2401
rect -903 -2435 -835 -2401
rect -745 -2435 -677 -2401
rect -587 -2435 -519 -2401
rect -429 -2435 -361 -2401
rect -271 -2435 -203 -2401
rect -113 -2435 -45 -2401
rect 45 -2435 113 -2401
rect 203 -2435 271 -2401
rect 361 -2435 429 -2401
rect 519 -2435 587 -2401
rect 677 -2435 745 -2401
rect 835 -2435 903 -2401
rect 993 -2435 1061 -2401
rect 1151 -2435 1219 -2401
<< metal1 >>
rect -1231 2435 -1139 2441
rect -1231 2401 -1219 2435
rect -1151 2401 -1139 2435
rect -1231 2395 -1139 2401
rect -1073 2435 -981 2441
rect -1073 2401 -1061 2435
rect -993 2401 -981 2435
rect -1073 2395 -981 2401
rect -915 2435 -823 2441
rect -915 2401 -903 2435
rect -835 2401 -823 2435
rect -915 2395 -823 2401
rect -757 2435 -665 2441
rect -757 2401 -745 2435
rect -677 2401 -665 2435
rect -757 2395 -665 2401
rect -599 2435 -507 2441
rect -599 2401 -587 2435
rect -519 2401 -507 2435
rect -599 2395 -507 2401
rect -441 2435 -349 2441
rect -441 2401 -429 2435
rect -361 2401 -349 2435
rect -441 2395 -349 2401
rect -283 2435 -191 2441
rect -283 2401 -271 2435
rect -203 2401 -191 2435
rect -283 2395 -191 2401
rect -125 2435 -33 2441
rect -125 2401 -113 2435
rect -45 2401 -33 2435
rect -125 2395 -33 2401
rect 33 2435 125 2441
rect 33 2401 45 2435
rect 113 2401 125 2435
rect 33 2395 125 2401
rect 191 2435 283 2441
rect 191 2401 203 2435
rect 271 2401 283 2435
rect 191 2395 283 2401
rect 349 2435 441 2441
rect 349 2401 361 2435
rect 429 2401 441 2435
rect 349 2395 441 2401
rect 507 2435 599 2441
rect 507 2401 519 2435
rect 587 2401 599 2435
rect 507 2395 599 2401
rect 665 2435 757 2441
rect 665 2401 677 2435
rect 745 2401 757 2435
rect 665 2395 757 2401
rect 823 2435 915 2441
rect 823 2401 835 2435
rect 903 2401 915 2435
rect 823 2395 915 2401
rect 981 2435 1073 2441
rect 981 2401 993 2435
rect 1061 2401 1073 2435
rect 981 2395 1073 2401
rect 1139 2435 1231 2441
rect 1139 2401 1151 2435
rect 1219 2401 1231 2435
rect 1139 2395 1231 2401
rect -1287 2351 -1241 2363
rect -1287 1975 -1281 2351
rect -1247 1975 -1241 2351
rect -1287 1963 -1241 1975
rect -1129 2351 -1083 2363
rect -1129 1975 -1123 2351
rect -1089 1975 -1083 2351
rect -1129 1963 -1083 1975
rect -971 2351 -925 2363
rect -971 1975 -965 2351
rect -931 1975 -925 2351
rect -971 1963 -925 1975
rect -813 2351 -767 2363
rect -813 1975 -807 2351
rect -773 1975 -767 2351
rect -813 1963 -767 1975
rect -655 2351 -609 2363
rect -655 1975 -649 2351
rect -615 1975 -609 2351
rect -655 1963 -609 1975
rect -497 2351 -451 2363
rect -497 1975 -491 2351
rect -457 1975 -451 2351
rect -497 1963 -451 1975
rect -339 2351 -293 2363
rect -339 1975 -333 2351
rect -299 1975 -293 2351
rect -339 1963 -293 1975
rect -181 2351 -135 2363
rect -181 1975 -175 2351
rect -141 1975 -135 2351
rect -181 1963 -135 1975
rect -23 2351 23 2363
rect -23 1975 -17 2351
rect 17 1975 23 2351
rect -23 1963 23 1975
rect 135 2351 181 2363
rect 135 1975 141 2351
rect 175 1975 181 2351
rect 135 1963 181 1975
rect 293 2351 339 2363
rect 293 1975 299 2351
rect 333 1975 339 2351
rect 293 1963 339 1975
rect 451 2351 497 2363
rect 451 1975 457 2351
rect 491 1975 497 2351
rect 451 1963 497 1975
rect 609 2351 655 2363
rect 609 1975 615 2351
rect 649 1975 655 2351
rect 609 1963 655 1975
rect 767 2351 813 2363
rect 767 1975 773 2351
rect 807 1975 813 2351
rect 767 1963 813 1975
rect 925 2351 971 2363
rect 925 1975 931 2351
rect 965 1975 971 2351
rect 925 1963 971 1975
rect 1083 2351 1129 2363
rect 1083 1975 1089 2351
rect 1123 1975 1129 2351
rect 1083 1963 1129 1975
rect 1241 2351 1287 2363
rect 1241 1975 1247 2351
rect 1281 1975 1287 2351
rect 1241 1963 1287 1975
rect -1231 1925 -1139 1931
rect -1231 1891 -1219 1925
rect -1151 1891 -1139 1925
rect -1231 1885 -1139 1891
rect -1073 1925 -981 1931
rect -1073 1891 -1061 1925
rect -993 1891 -981 1925
rect -1073 1885 -981 1891
rect -915 1925 -823 1931
rect -915 1891 -903 1925
rect -835 1891 -823 1925
rect -915 1885 -823 1891
rect -757 1925 -665 1931
rect -757 1891 -745 1925
rect -677 1891 -665 1925
rect -757 1885 -665 1891
rect -599 1925 -507 1931
rect -599 1891 -587 1925
rect -519 1891 -507 1925
rect -599 1885 -507 1891
rect -441 1925 -349 1931
rect -441 1891 -429 1925
rect -361 1891 -349 1925
rect -441 1885 -349 1891
rect -283 1925 -191 1931
rect -283 1891 -271 1925
rect -203 1891 -191 1925
rect -283 1885 -191 1891
rect -125 1925 -33 1931
rect -125 1891 -113 1925
rect -45 1891 -33 1925
rect -125 1885 -33 1891
rect 33 1925 125 1931
rect 33 1891 45 1925
rect 113 1891 125 1925
rect 33 1885 125 1891
rect 191 1925 283 1931
rect 191 1891 203 1925
rect 271 1891 283 1925
rect 191 1885 283 1891
rect 349 1925 441 1931
rect 349 1891 361 1925
rect 429 1891 441 1925
rect 349 1885 441 1891
rect 507 1925 599 1931
rect 507 1891 519 1925
rect 587 1891 599 1925
rect 507 1885 599 1891
rect 665 1925 757 1931
rect 665 1891 677 1925
rect 745 1891 757 1925
rect 665 1885 757 1891
rect 823 1925 915 1931
rect 823 1891 835 1925
rect 903 1891 915 1925
rect 823 1885 915 1891
rect 981 1925 1073 1931
rect 981 1891 993 1925
rect 1061 1891 1073 1925
rect 981 1885 1073 1891
rect 1139 1925 1231 1931
rect 1139 1891 1151 1925
rect 1219 1891 1231 1925
rect 1139 1885 1231 1891
rect -1231 1817 -1139 1823
rect -1231 1783 -1219 1817
rect -1151 1783 -1139 1817
rect -1231 1777 -1139 1783
rect -1073 1817 -981 1823
rect -1073 1783 -1061 1817
rect -993 1783 -981 1817
rect -1073 1777 -981 1783
rect -915 1817 -823 1823
rect -915 1783 -903 1817
rect -835 1783 -823 1817
rect -915 1777 -823 1783
rect -757 1817 -665 1823
rect -757 1783 -745 1817
rect -677 1783 -665 1817
rect -757 1777 -665 1783
rect -599 1817 -507 1823
rect -599 1783 -587 1817
rect -519 1783 -507 1817
rect -599 1777 -507 1783
rect -441 1817 -349 1823
rect -441 1783 -429 1817
rect -361 1783 -349 1817
rect -441 1777 -349 1783
rect -283 1817 -191 1823
rect -283 1783 -271 1817
rect -203 1783 -191 1817
rect -283 1777 -191 1783
rect -125 1817 -33 1823
rect -125 1783 -113 1817
rect -45 1783 -33 1817
rect -125 1777 -33 1783
rect 33 1817 125 1823
rect 33 1783 45 1817
rect 113 1783 125 1817
rect 33 1777 125 1783
rect 191 1817 283 1823
rect 191 1783 203 1817
rect 271 1783 283 1817
rect 191 1777 283 1783
rect 349 1817 441 1823
rect 349 1783 361 1817
rect 429 1783 441 1817
rect 349 1777 441 1783
rect 507 1817 599 1823
rect 507 1783 519 1817
rect 587 1783 599 1817
rect 507 1777 599 1783
rect 665 1817 757 1823
rect 665 1783 677 1817
rect 745 1783 757 1817
rect 665 1777 757 1783
rect 823 1817 915 1823
rect 823 1783 835 1817
rect 903 1783 915 1817
rect 823 1777 915 1783
rect 981 1817 1073 1823
rect 981 1783 993 1817
rect 1061 1783 1073 1817
rect 981 1777 1073 1783
rect 1139 1817 1231 1823
rect 1139 1783 1151 1817
rect 1219 1783 1231 1817
rect 1139 1777 1231 1783
rect -1287 1733 -1241 1745
rect -1287 1357 -1281 1733
rect -1247 1357 -1241 1733
rect -1287 1345 -1241 1357
rect -1129 1733 -1083 1745
rect -1129 1357 -1123 1733
rect -1089 1357 -1083 1733
rect -1129 1345 -1083 1357
rect -971 1733 -925 1745
rect -971 1357 -965 1733
rect -931 1357 -925 1733
rect -971 1345 -925 1357
rect -813 1733 -767 1745
rect -813 1357 -807 1733
rect -773 1357 -767 1733
rect -813 1345 -767 1357
rect -655 1733 -609 1745
rect -655 1357 -649 1733
rect -615 1357 -609 1733
rect -655 1345 -609 1357
rect -497 1733 -451 1745
rect -497 1357 -491 1733
rect -457 1357 -451 1733
rect -497 1345 -451 1357
rect -339 1733 -293 1745
rect -339 1357 -333 1733
rect -299 1357 -293 1733
rect -339 1345 -293 1357
rect -181 1733 -135 1745
rect -181 1357 -175 1733
rect -141 1357 -135 1733
rect -181 1345 -135 1357
rect -23 1733 23 1745
rect -23 1357 -17 1733
rect 17 1357 23 1733
rect -23 1345 23 1357
rect 135 1733 181 1745
rect 135 1357 141 1733
rect 175 1357 181 1733
rect 135 1345 181 1357
rect 293 1733 339 1745
rect 293 1357 299 1733
rect 333 1357 339 1733
rect 293 1345 339 1357
rect 451 1733 497 1745
rect 451 1357 457 1733
rect 491 1357 497 1733
rect 451 1345 497 1357
rect 609 1733 655 1745
rect 609 1357 615 1733
rect 649 1357 655 1733
rect 609 1345 655 1357
rect 767 1733 813 1745
rect 767 1357 773 1733
rect 807 1357 813 1733
rect 767 1345 813 1357
rect 925 1733 971 1745
rect 925 1357 931 1733
rect 965 1357 971 1733
rect 925 1345 971 1357
rect 1083 1733 1129 1745
rect 1083 1357 1089 1733
rect 1123 1357 1129 1733
rect 1083 1345 1129 1357
rect 1241 1733 1287 1745
rect 1241 1357 1247 1733
rect 1281 1357 1287 1733
rect 1241 1345 1287 1357
rect -1231 1307 -1139 1313
rect -1231 1273 -1219 1307
rect -1151 1273 -1139 1307
rect -1231 1267 -1139 1273
rect -1073 1307 -981 1313
rect -1073 1273 -1061 1307
rect -993 1273 -981 1307
rect -1073 1267 -981 1273
rect -915 1307 -823 1313
rect -915 1273 -903 1307
rect -835 1273 -823 1307
rect -915 1267 -823 1273
rect -757 1307 -665 1313
rect -757 1273 -745 1307
rect -677 1273 -665 1307
rect -757 1267 -665 1273
rect -599 1307 -507 1313
rect -599 1273 -587 1307
rect -519 1273 -507 1307
rect -599 1267 -507 1273
rect -441 1307 -349 1313
rect -441 1273 -429 1307
rect -361 1273 -349 1307
rect -441 1267 -349 1273
rect -283 1307 -191 1313
rect -283 1273 -271 1307
rect -203 1273 -191 1307
rect -283 1267 -191 1273
rect -125 1307 -33 1313
rect -125 1273 -113 1307
rect -45 1273 -33 1307
rect -125 1267 -33 1273
rect 33 1307 125 1313
rect 33 1273 45 1307
rect 113 1273 125 1307
rect 33 1267 125 1273
rect 191 1307 283 1313
rect 191 1273 203 1307
rect 271 1273 283 1307
rect 191 1267 283 1273
rect 349 1307 441 1313
rect 349 1273 361 1307
rect 429 1273 441 1307
rect 349 1267 441 1273
rect 507 1307 599 1313
rect 507 1273 519 1307
rect 587 1273 599 1307
rect 507 1267 599 1273
rect 665 1307 757 1313
rect 665 1273 677 1307
rect 745 1273 757 1307
rect 665 1267 757 1273
rect 823 1307 915 1313
rect 823 1273 835 1307
rect 903 1273 915 1307
rect 823 1267 915 1273
rect 981 1307 1073 1313
rect 981 1273 993 1307
rect 1061 1273 1073 1307
rect 981 1267 1073 1273
rect 1139 1307 1231 1313
rect 1139 1273 1151 1307
rect 1219 1273 1231 1307
rect 1139 1267 1231 1273
rect -1231 1199 -1139 1205
rect -1231 1165 -1219 1199
rect -1151 1165 -1139 1199
rect -1231 1159 -1139 1165
rect -1073 1199 -981 1205
rect -1073 1165 -1061 1199
rect -993 1165 -981 1199
rect -1073 1159 -981 1165
rect -915 1199 -823 1205
rect -915 1165 -903 1199
rect -835 1165 -823 1199
rect -915 1159 -823 1165
rect -757 1199 -665 1205
rect -757 1165 -745 1199
rect -677 1165 -665 1199
rect -757 1159 -665 1165
rect -599 1199 -507 1205
rect -599 1165 -587 1199
rect -519 1165 -507 1199
rect -599 1159 -507 1165
rect -441 1199 -349 1205
rect -441 1165 -429 1199
rect -361 1165 -349 1199
rect -441 1159 -349 1165
rect -283 1199 -191 1205
rect -283 1165 -271 1199
rect -203 1165 -191 1199
rect -283 1159 -191 1165
rect -125 1199 -33 1205
rect -125 1165 -113 1199
rect -45 1165 -33 1199
rect -125 1159 -33 1165
rect 33 1199 125 1205
rect 33 1165 45 1199
rect 113 1165 125 1199
rect 33 1159 125 1165
rect 191 1199 283 1205
rect 191 1165 203 1199
rect 271 1165 283 1199
rect 191 1159 283 1165
rect 349 1199 441 1205
rect 349 1165 361 1199
rect 429 1165 441 1199
rect 349 1159 441 1165
rect 507 1199 599 1205
rect 507 1165 519 1199
rect 587 1165 599 1199
rect 507 1159 599 1165
rect 665 1199 757 1205
rect 665 1165 677 1199
rect 745 1165 757 1199
rect 665 1159 757 1165
rect 823 1199 915 1205
rect 823 1165 835 1199
rect 903 1165 915 1199
rect 823 1159 915 1165
rect 981 1199 1073 1205
rect 981 1165 993 1199
rect 1061 1165 1073 1199
rect 981 1159 1073 1165
rect 1139 1199 1231 1205
rect 1139 1165 1151 1199
rect 1219 1165 1231 1199
rect 1139 1159 1231 1165
rect -1287 1115 -1241 1127
rect -1287 739 -1281 1115
rect -1247 739 -1241 1115
rect -1287 727 -1241 739
rect -1129 1115 -1083 1127
rect -1129 739 -1123 1115
rect -1089 739 -1083 1115
rect -1129 727 -1083 739
rect -971 1115 -925 1127
rect -971 739 -965 1115
rect -931 739 -925 1115
rect -971 727 -925 739
rect -813 1115 -767 1127
rect -813 739 -807 1115
rect -773 739 -767 1115
rect -813 727 -767 739
rect -655 1115 -609 1127
rect -655 739 -649 1115
rect -615 739 -609 1115
rect -655 727 -609 739
rect -497 1115 -451 1127
rect -497 739 -491 1115
rect -457 739 -451 1115
rect -497 727 -451 739
rect -339 1115 -293 1127
rect -339 739 -333 1115
rect -299 739 -293 1115
rect -339 727 -293 739
rect -181 1115 -135 1127
rect -181 739 -175 1115
rect -141 739 -135 1115
rect -181 727 -135 739
rect -23 1115 23 1127
rect -23 739 -17 1115
rect 17 739 23 1115
rect -23 727 23 739
rect 135 1115 181 1127
rect 135 739 141 1115
rect 175 739 181 1115
rect 135 727 181 739
rect 293 1115 339 1127
rect 293 739 299 1115
rect 333 739 339 1115
rect 293 727 339 739
rect 451 1115 497 1127
rect 451 739 457 1115
rect 491 739 497 1115
rect 451 727 497 739
rect 609 1115 655 1127
rect 609 739 615 1115
rect 649 739 655 1115
rect 609 727 655 739
rect 767 1115 813 1127
rect 767 739 773 1115
rect 807 739 813 1115
rect 767 727 813 739
rect 925 1115 971 1127
rect 925 739 931 1115
rect 965 739 971 1115
rect 925 727 971 739
rect 1083 1115 1129 1127
rect 1083 739 1089 1115
rect 1123 739 1129 1115
rect 1083 727 1129 739
rect 1241 1115 1287 1127
rect 1241 739 1247 1115
rect 1281 739 1287 1115
rect 1241 727 1287 739
rect -1231 689 -1139 695
rect -1231 655 -1219 689
rect -1151 655 -1139 689
rect -1231 649 -1139 655
rect -1073 689 -981 695
rect -1073 655 -1061 689
rect -993 655 -981 689
rect -1073 649 -981 655
rect -915 689 -823 695
rect -915 655 -903 689
rect -835 655 -823 689
rect -915 649 -823 655
rect -757 689 -665 695
rect -757 655 -745 689
rect -677 655 -665 689
rect -757 649 -665 655
rect -599 689 -507 695
rect -599 655 -587 689
rect -519 655 -507 689
rect -599 649 -507 655
rect -441 689 -349 695
rect -441 655 -429 689
rect -361 655 -349 689
rect -441 649 -349 655
rect -283 689 -191 695
rect -283 655 -271 689
rect -203 655 -191 689
rect -283 649 -191 655
rect -125 689 -33 695
rect -125 655 -113 689
rect -45 655 -33 689
rect -125 649 -33 655
rect 33 689 125 695
rect 33 655 45 689
rect 113 655 125 689
rect 33 649 125 655
rect 191 689 283 695
rect 191 655 203 689
rect 271 655 283 689
rect 191 649 283 655
rect 349 689 441 695
rect 349 655 361 689
rect 429 655 441 689
rect 349 649 441 655
rect 507 689 599 695
rect 507 655 519 689
rect 587 655 599 689
rect 507 649 599 655
rect 665 689 757 695
rect 665 655 677 689
rect 745 655 757 689
rect 665 649 757 655
rect 823 689 915 695
rect 823 655 835 689
rect 903 655 915 689
rect 823 649 915 655
rect 981 689 1073 695
rect 981 655 993 689
rect 1061 655 1073 689
rect 981 649 1073 655
rect 1139 689 1231 695
rect 1139 655 1151 689
rect 1219 655 1231 689
rect 1139 649 1231 655
rect -1231 581 -1139 587
rect -1231 547 -1219 581
rect -1151 547 -1139 581
rect -1231 541 -1139 547
rect -1073 581 -981 587
rect -1073 547 -1061 581
rect -993 547 -981 581
rect -1073 541 -981 547
rect -915 581 -823 587
rect -915 547 -903 581
rect -835 547 -823 581
rect -915 541 -823 547
rect -757 581 -665 587
rect -757 547 -745 581
rect -677 547 -665 581
rect -757 541 -665 547
rect -599 581 -507 587
rect -599 547 -587 581
rect -519 547 -507 581
rect -599 541 -507 547
rect -441 581 -349 587
rect -441 547 -429 581
rect -361 547 -349 581
rect -441 541 -349 547
rect -283 581 -191 587
rect -283 547 -271 581
rect -203 547 -191 581
rect -283 541 -191 547
rect -125 581 -33 587
rect -125 547 -113 581
rect -45 547 -33 581
rect -125 541 -33 547
rect 33 581 125 587
rect 33 547 45 581
rect 113 547 125 581
rect 33 541 125 547
rect 191 581 283 587
rect 191 547 203 581
rect 271 547 283 581
rect 191 541 283 547
rect 349 581 441 587
rect 349 547 361 581
rect 429 547 441 581
rect 349 541 441 547
rect 507 581 599 587
rect 507 547 519 581
rect 587 547 599 581
rect 507 541 599 547
rect 665 581 757 587
rect 665 547 677 581
rect 745 547 757 581
rect 665 541 757 547
rect 823 581 915 587
rect 823 547 835 581
rect 903 547 915 581
rect 823 541 915 547
rect 981 581 1073 587
rect 981 547 993 581
rect 1061 547 1073 581
rect 981 541 1073 547
rect 1139 581 1231 587
rect 1139 547 1151 581
rect 1219 547 1231 581
rect 1139 541 1231 547
rect -1287 497 -1241 509
rect -1287 121 -1281 497
rect -1247 121 -1241 497
rect -1287 109 -1241 121
rect -1129 497 -1083 509
rect -1129 121 -1123 497
rect -1089 121 -1083 497
rect -1129 109 -1083 121
rect -971 497 -925 509
rect -971 121 -965 497
rect -931 121 -925 497
rect -971 109 -925 121
rect -813 497 -767 509
rect -813 121 -807 497
rect -773 121 -767 497
rect -813 109 -767 121
rect -655 497 -609 509
rect -655 121 -649 497
rect -615 121 -609 497
rect -655 109 -609 121
rect -497 497 -451 509
rect -497 121 -491 497
rect -457 121 -451 497
rect -497 109 -451 121
rect -339 497 -293 509
rect -339 121 -333 497
rect -299 121 -293 497
rect -339 109 -293 121
rect -181 497 -135 509
rect -181 121 -175 497
rect -141 121 -135 497
rect -181 109 -135 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 135 497 181 509
rect 135 121 141 497
rect 175 121 181 497
rect 135 109 181 121
rect 293 497 339 509
rect 293 121 299 497
rect 333 121 339 497
rect 293 109 339 121
rect 451 497 497 509
rect 451 121 457 497
rect 491 121 497 497
rect 451 109 497 121
rect 609 497 655 509
rect 609 121 615 497
rect 649 121 655 497
rect 609 109 655 121
rect 767 497 813 509
rect 767 121 773 497
rect 807 121 813 497
rect 767 109 813 121
rect 925 497 971 509
rect 925 121 931 497
rect 965 121 971 497
rect 925 109 971 121
rect 1083 497 1129 509
rect 1083 121 1089 497
rect 1123 121 1129 497
rect 1083 109 1129 121
rect 1241 497 1287 509
rect 1241 121 1247 497
rect 1281 121 1287 497
rect 1241 109 1287 121
rect -1231 71 -1139 77
rect -1231 37 -1219 71
rect -1151 37 -1139 71
rect -1231 31 -1139 37
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect 1139 71 1231 77
rect 1139 37 1151 71
rect 1219 37 1231 71
rect 1139 31 1231 37
rect -1231 -37 -1139 -31
rect -1231 -71 -1219 -37
rect -1151 -71 -1139 -37
rect -1231 -77 -1139 -71
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect 1139 -37 1231 -31
rect 1139 -71 1151 -37
rect 1219 -71 1231 -37
rect 1139 -77 1231 -71
rect -1287 -121 -1241 -109
rect -1287 -497 -1281 -121
rect -1247 -497 -1241 -121
rect -1287 -509 -1241 -497
rect -1129 -121 -1083 -109
rect -1129 -497 -1123 -121
rect -1089 -497 -1083 -121
rect -1129 -509 -1083 -497
rect -971 -121 -925 -109
rect -971 -497 -965 -121
rect -931 -497 -925 -121
rect -971 -509 -925 -497
rect -813 -121 -767 -109
rect -813 -497 -807 -121
rect -773 -497 -767 -121
rect -813 -509 -767 -497
rect -655 -121 -609 -109
rect -655 -497 -649 -121
rect -615 -497 -609 -121
rect -655 -509 -609 -497
rect -497 -121 -451 -109
rect -497 -497 -491 -121
rect -457 -497 -451 -121
rect -497 -509 -451 -497
rect -339 -121 -293 -109
rect -339 -497 -333 -121
rect -299 -497 -293 -121
rect -339 -509 -293 -497
rect -181 -121 -135 -109
rect -181 -497 -175 -121
rect -141 -497 -135 -121
rect -181 -509 -135 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 135 -121 181 -109
rect 135 -497 141 -121
rect 175 -497 181 -121
rect 135 -509 181 -497
rect 293 -121 339 -109
rect 293 -497 299 -121
rect 333 -497 339 -121
rect 293 -509 339 -497
rect 451 -121 497 -109
rect 451 -497 457 -121
rect 491 -497 497 -121
rect 451 -509 497 -497
rect 609 -121 655 -109
rect 609 -497 615 -121
rect 649 -497 655 -121
rect 609 -509 655 -497
rect 767 -121 813 -109
rect 767 -497 773 -121
rect 807 -497 813 -121
rect 767 -509 813 -497
rect 925 -121 971 -109
rect 925 -497 931 -121
rect 965 -497 971 -121
rect 925 -509 971 -497
rect 1083 -121 1129 -109
rect 1083 -497 1089 -121
rect 1123 -497 1129 -121
rect 1083 -509 1129 -497
rect 1241 -121 1287 -109
rect 1241 -497 1247 -121
rect 1281 -497 1287 -121
rect 1241 -509 1287 -497
rect -1231 -547 -1139 -541
rect -1231 -581 -1219 -547
rect -1151 -581 -1139 -547
rect -1231 -587 -1139 -581
rect -1073 -547 -981 -541
rect -1073 -581 -1061 -547
rect -993 -581 -981 -547
rect -1073 -587 -981 -581
rect -915 -547 -823 -541
rect -915 -581 -903 -547
rect -835 -581 -823 -547
rect -915 -587 -823 -581
rect -757 -547 -665 -541
rect -757 -581 -745 -547
rect -677 -581 -665 -547
rect -757 -587 -665 -581
rect -599 -547 -507 -541
rect -599 -581 -587 -547
rect -519 -581 -507 -547
rect -599 -587 -507 -581
rect -441 -547 -349 -541
rect -441 -581 -429 -547
rect -361 -581 -349 -547
rect -441 -587 -349 -581
rect -283 -547 -191 -541
rect -283 -581 -271 -547
rect -203 -581 -191 -547
rect -283 -587 -191 -581
rect -125 -547 -33 -541
rect -125 -581 -113 -547
rect -45 -581 -33 -547
rect -125 -587 -33 -581
rect 33 -547 125 -541
rect 33 -581 45 -547
rect 113 -581 125 -547
rect 33 -587 125 -581
rect 191 -547 283 -541
rect 191 -581 203 -547
rect 271 -581 283 -547
rect 191 -587 283 -581
rect 349 -547 441 -541
rect 349 -581 361 -547
rect 429 -581 441 -547
rect 349 -587 441 -581
rect 507 -547 599 -541
rect 507 -581 519 -547
rect 587 -581 599 -547
rect 507 -587 599 -581
rect 665 -547 757 -541
rect 665 -581 677 -547
rect 745 -581 757 -547
rect 665 -587 757 -581
rect 823 -547 915 -541
rect 823 -581 835 -547
rect 903 -581 915 -547
rect 823 -587 915 -581
rect 981 -547 1073 -541
rect 981 -581 993 -547
rect 1061 -581 1073 -547
rect 981 -587 1073 -581
rect 1139 -547 1231 -541
rect 1139 -581 1151 -547
rect 1219 -581 1231 -547
rect 1139 -587 1231 -581
rect -1231 -655 -1139 -649
rect -1231 -689 -1219 -655
rect -1151 -689 -1139 -655
rect -1231 -695 -1139 -689
rect -1073 -655 -981 -649
rect -1073 -689 -1061 -655
rect -993 -689 -981 -655
rect -1073 -695 -981 -689
rect -915 -655 -823 -649
rect -915 -689 -903 -655
rect -835 -689 -823 -655
rect -915 -695 -823 -689
rect -757 -655 -665 -649
rect -757 -689 -745 -655
rect -677 -689 -665 -655
rect -757 -695 -665 -689
rect -599 -655 -507 -649
rect -599 -689 -587 -655
rect -519 -689 -507 -655
rect -599 -695 -507 -689
rect -441 -655 -349 -649
rect -441 -689 -429 -655
rect -361 -689 -349 -655
rect -441 -695 -349 -689
rect -283 -655 -191 -649
rect -283 -689 -271 -655
rect -203 -689 -191 -655
rect -283 -695 -191 -689
rect -125 -655 -33 -649
rect -125 -689 -113 -655
rect -45 -689 -33 -655
rect -125 -695 -33 -689
rect 33 -655 125 -649
rect 33 -689 45 -655
rect 113 -689 125 -655
rect 33 -695 125 -689
rect 191 -655 283 -649
rect 191 -689 203 -655
rect 271 -689 283 -655
rect 191 -695 283 -689
rect 349 -655 441 -649
rect 349 -689 361 -655
rect 429 -689 441 -655
rect 349 -695 441 -689
rect 507 -655 599 -649
rect 507 -689 519 -655
rect 587 -689 599 -655
rect 507 -695 599 -689
rect 665 -655 757 -649
rect 665 -689 677 -655
rect 745 -689 757 -655
rect 665 -695 757 -689
rect 823 -655 915 -649
rect 823 -689 835 -655
rect 903 -689 915 -655
rect 823 -695 915 -689
rect 981 -655 1073 -649
rect 981 -689 993 -655
rect 1061 -689 1073 -655
rect 981 -695 1073 -689
rect 1139 -655 1231 -649
rect 1139 -689 1151 -655
rect 1219 -689 1231 -655
rect 1139 -695 1231 -689
rect -1287 -739 -1241 -727
rect -1287 -1115 -1281 -739
rect -1247 -1115 -1241 -739
rect -1287 -1127 -1241 -1115
rect -1129 -739 -1083 -727
rect -1129 -1115 -1123 -739
rect -1089 -1115 -1083 -739
rect -1129 -1127 -1083 -1115
rect -971 -739 -925 -727
rect -971 -1115 -965 -739
rect -931 -1115 -925 -739
rect -971 -1127 -925 -1115
rect -813 -739 -767 -727
rect -813 -1115 -807 -739
rect -773 -1115 -767 -739
rect -813 -1127 -767 -1115
rect -655 -739 -609 -727
rect -655 -1115 -649 -739
rect -615 -1115 -609 -739
rect -655 -1127 -609 -1115
rect -497 -739 -451 -727
rect -497 -1115 -491 -739
rect -457 -1115 -451 -739
rect -497 -1127 -451 -1115
rect -339 -739 -293 -727
rect -339 -1115 -333 -739
rect -299 -1115 -293 -739
rect -339 -1127 -293 -1115
rect -181 -739 -135 -727
rect -181 -1115 -175 -739
rect -141 -1115 -135 -739
rect -181 -1127 -135 -1115
rect -23 -739 23 -727
rect -23 -1115 -17 -739
rect 17 -1115 23 -739
rect -23 -1127 23 -1115
rect 135 -739 181 -727
rect 135 -1115 141 -739
rect 175 -1115 181 -739
rect 135 -1127 181 -1115
rect 293 -739 339 -727
rect 293 -1115 299 -739
rect 333 -1115 339 -739
rect 293 -1127 339 -1115
rect 451 -739 497 -727
rect 451 -1115 457 -739
rect 491 -1115 497 -739
rect 451 -1127 497 -1115
rect 609 -739 655 -727
rect 609 -1115 615 -739
rect 649 -1115 655 -739
rect 609 -1127 655 -1115
rect 767 -739 813 -727
rect 767 -1115 773 -739
rect 807 -1115 813 -739
rect 767 -1127 813 -1115
rect 925 -739 971 -727
rect 925 -1115 931 -739
rect 965 -1115 971 -739
rect 925 -1127 971 -1115
rect 1083 -739 1129 -727
rect 1083 -1115 1089 -739
rect 1123 -1115 1129 -739
rect 1083 -1127 1129 -1115
rect 1241 -739 1287 -727
rect 1241 -1115 1247 -739
rect 1281 -1115 1287 -739
rect 1241 -1127 1287 -1115
rect -1231 -1165 -1139 -1159
rect -1231 -1199 -1219 -1165
rect -1151 -1199 -1139 -1165
rect -1231 -1205 -1139 -1199
rect -1073 -1165 -981 -1159
rect -1073 -1199 -1061 -1165
rect -993 -1199 -981 -1165
rect -1073 -1205 -981 -1199
rect -915 -1165 -823 -1159
rect -915 -1199 -903 -1165
rect -835 -1199 -823 -1165
rect -915 -1205 -823 -1199
rect -757 -1165 -665 -1159
rect -757 -1199 -745 -1165
rect -677 -1199 -665 -1165
rect -757 -1205 -665 -1199
rect -599 -1165 -507 -1159
rect -599 -1199 -587 -1165
rect -519 -1199 -507 -1165
rect -599 -1205 -507 -1199
rect -441 -1165 -349 -1159
rect -441 -1199 -429 -1165
rect -361 -1199 -349 -1165
rect -441 -1205 -349 -1199
rect -283 -1165 -191 -1159
rect -283 -1199 -271 -1165
rect -203 -1199 -191 -1165
rect -283 -1205 -191 -1199
rect -125 -1165 -33 -1159
rect -125 -1199 -113 -1165
rect -45 -1199 -33 -1165
rect -125 -1205 -33 -1199
rect 33 -1165 125 -1159
rect 33 -1199 45 -1165
rect 113 -1199 125 -1165
rect 33 -1205 125 -1199
rect 191 -1165 283 -1159
rect 191 -1199 203 -1165
rect 271 -1199 283 -1165
rect 191 -1205 283 -1199
rect 349 -1165 441 -1159
rect 349 -1199 361 -1165
rect 429 -1199 441 -1165
rect 349 -1205 441 -1199
rect 507 -1165 599 -1159
rect 507 -1199 519 -1165
rect 587 -1199 599 -1165
rect 507 -1205 599 -1199
rect 665 -1165 757 -1159
rect 665 -1199 677 -1165
rect 745 -1199 757 -1165
rect 665 -1205 757 -1199
rect 823 -1165 915 -1159
rect 823 -1199 835 -1165
rect 903 -1199 915 -1165
rect 823 -1205 915 -1199
rect 981 -1165 1073 -1159
rect 981 -1199 993 -1165
rect 1061 -1199 1073 -1165
rect 981 -1205 1073 -1199
rect 1139 -1165 1231 -1159
rect 1139 -1199 1151 -1165
rect 1219 -1199 1231 -1165
rect 1139 -1205 1231 -1199
rect -1231 -1273 -1139 -1267
rect -1231 -1307 -1219 -1273
rect -1151 -1307 -1139 -1273
rect -1231 -1313 -1139 -1307
rect -1073 -1273 -981 -1267
rect -1073 -1307 -1061 -1273
rect -993 -1307 -981 -1273
rect -1073 -1313 -981 -1307
rect -915 -1273 -823 -1267
rect -915 -1307 -903 -1273
rect -835 -1307 -823 -1273
rect -915 -1313 -823 -1307
rect -757 -1273 -665 -1267
rect -757 -1307 -745 -1273
rect -677 -1307 -665 -1273
rect -757 -1313 -665 -1307
rect -599 -1273 -507 -1267
rect -599 -1307 -587 -1273
rect -519 -1307 -507 -1273
rect -599 -1313 -507 -1307
rect -441 -1273 -349 -1267
rect -441 -1307 -429 -1273
rect -361 -1307 -349 -1273
rect -441 -1313 -349 -1307
rect -283 -1273 -191 -1267
rect -283 -1307 -271 -1273
rect -203 -1307 -191 -1273
rect -283 -1313 -191 -1307
rect -125 -1273 -33 -1267
rect -125 -1307 -113 -1273
rect -45 -1307 -33 -1273
rect -125 -1313 -33 -1307
rect 33 -1273 125 -1267
rect 33 -1307 45 -1273
rect 113 -1307 125 -1273
rect 33 -1313 125 -1307
rect 191 -1273 283 -1267
rect 191 -1307 203 -1273
rect 271 -1307 283 -1273
rect 191 -1313 283 -1307
rect 349 -1273 441 -1267
rect 349 -1307 361 -1273
rect 429 -1307 441 -1273
rect 349 -1313 441 -1307
rect 507 -1273 599 -1267
rect 507 -1307 519 -1273
rect 587 -1307 599 -1273
rect 507 -1313 599 -1307
rect 665 -1273 757 -1267
rect 665 -1307 677 -1273
rect 745 -1307 757 -1273
rect 665 -1313 757 -1307
rect 823 -1273 915 -1267
rect 823 -1307 835 -1273
rect 903 -1307 915 -1273
rect 823 -1313 915 -1307
rect 981 -1273 1073 -1267
rect 981 -1307 993 -1273
rect 1061 -1307 1073 -1273
rect 981 -1313 1073 -1307
rect 1139 -1273 1231 -1267
rect 1139 -1307 1151 -1273
rect 1219 -1307 1231 -1273
rect 1139 -1313 1231 -1307
rect -1287 -1357 -1241 -1345
rect -1287 -1733 -1281 -1357
rect -1247 -1733 -1241 -1357
rect -1287 -1745 -1241 -1733
rect -1129 -1357 -1083 -1345
rect -1129 -1733 -1123 -1357
rect -1089 -1733 -1083 -1357
rect -1129 -1745 -1083 -1733
rect -971 -1357 -925 -1345
rect -971 -1733 -965 -1357
rect -931 -1733 -925 -1357
rect -971 -1745 -925 -1733
rect -813 -1357 -767 -1345
rect -813 -1733 -807 -1357
rect -773 -1733 -767 -1357
rect -813 -1745 -767 -1733
rect -655 -1357 -609 -1345
rect -655 -1733 -649 -1357
rect -615 -1733 -609 -1357
rect -655 -1745 -609 -1733
rect -497 -1357 -451 -1345
rect -497 -1733 -491 -1357
rect -457 -1733 -451 -1357
rect -497 -1745 -451 -1733
rect -339 -1357 -293 -1345
rect -339 -1733 -333 -1357
rect -299 -1733 -293 -1357
rect -339 -1745 -293 -1733
rect -181 -1357 -135 -1345
rect -181 -1733 -175 -1357
rect -141 -1733 -135 -1357
rect -181 -1745 -135 -1733
rect -23 -1357 23 -1345
rect -23 -1733 -17 -1357
rect 17 -1733 23 -1357
rect -23 -1745 23 -1733
rect 135 -1357 181 -1345
rect 135 -1733 141 -1357
rect 175 -1733 181 -1357
rect 135 -1745 181 -1733
rect 293 -1357 339 -1345
rect 293 -1733 299 -1357
rect 333 -1733 339 -1357
rect 293 -1745 339 -1733
rect 451 -1357 497 -1345
rect 451 -1733 457 -1357
rect 491 -1733 497 -1357
rect 451 -1745 497 -1733
rect 609 -1357 655 -1345
rect 609 -1733 615 -1357
rect 649 -1733 655 -1357
rect 609 -1745 655 -1733
rect 767 -1357 813 -1345
rect 767 -1733 773 -1357
rect 807 -1733 813 -1357
rect 767 -1745 813 -1733
rect 925 -1357 971 -1345
rect 925 -1733 931 -1357
rect 965 -1733 971 -1357
rect 925 -1745 971 -1733
rect 1083 -1357 1129 -1345
rect 1083 -1733 1089 -1357
rect 1123 -1733 1129 -1357
rect 1083 -1745 1129 -1733
rect 1241 -1357 1287 -1345
rect 1241 -1733 1247 -1357
rect 1281 -1733 1287 -1357
rect 1241 -1745 1287 -1733
rect -1231 -1783 -1139 -1777
rect -1231 -1817 -1219 -1783
rect -1151 -1817 -1139 -1783
rect -1231 -1823 -1139 -1817
rect -1073 -1783 -981 -1777
rect -1073 -1817 -1061 -1783
rect -993 -1817 -981 -1783
rect -1073 -1823 -981 -1817
rect -915 -1783 -823 -1777
rect -915 -1817 -903 -1783
rect -835 -1817 -823 -1783
rect -915 -1823 -823 -1817
rect -757 -1783 -665 -1777
rect -757 -1817 -745 -1783
rect -677 -1817 -665 -1783
rect -757 -1823 -665 -1817
rect -599 -1783 -507 -1777
rect -599 -1817 -587 -1783
rect -519 -1817 -507 -1783
rect -599 -1823 -507 -1817
rect -441 -1783 -349 -1777
rect -441 -1817 -429 -1783
rect -361 -1817 -349 -1783
rect -441 -1823 -349 -1817
rect -283 -1783 -191 -1777
rect -283 -1817 -271 -1783
rect -203 -1817 -191 -1783
rect -283 -1823 -191 -1817
rect -125 -1783 -33 -1777
rect -125 -1817 -113 -1783
rect -45 -1817 -33 -1783
rect -125 -1823 -33 -1817
rect 33 -1783 125 -1777
rect 33 -1817 45 -1783
rect 113 -1817 125 -1783
rect 33 -1823 125 -1817
rect 191 -1783 283 -1777
rect 191 -1817 203 -1783
rect 271 -1817 283 -1783
rect 191 -1823 283 -1817
rect 349 -1783 441 -1777
rect 349 -1817 361 -1783
rect 429 -1817 441 -1783
rect 349 -1823 441 -1817
rect 507 -1783 599 -1777
rect 507 -1817 519 -1783
rect 587 -1817 599 -1783
rect 507 -1823 599 -1817
rect 665 -1783 757 -1777
rect 665 -1817 677 -1783
rect 745 -1817 757 -1783
rect 665 -1823 757 -1817
rect 823 -1783 915 -1777
rect 823 -1817 835 -1783
rect 903 -1817 915 -1783
rect 823 -1823 915 -1817
rect 981 -1783 1073 -1777
rect 981 -1817 993 -1783
rect 1061 -1817 1073 -1783
rect 981 -1823 1073 -1817
rect 1139 -1783 1231 -1777
rect 1139 -1817 1151 -1783
rect 1219 -1817 1231 -1783
rect 1139 -1823 1231 -1817
rect -1231 -1891 -1139 -1885
rect -1231 -1925 -1219 -1891
rect -1151 -1925 -1139 -1891
rect -1231 -1931 -1139 -1925
rect -1073 -1891 -981 -1885
rect -1073 -1925 -1061 -1891
rect -993 -1925 -981 -1891
rect -1073 -1931 -981 -1925
rect -915 -1891 -823 -1885
rect -915 -1925 -903 -1891
rect -835 -1925 -823 -1891
rect -915 -1931 -823 -1925
rect -757 -1891 -665 -1885
rect -757 -1925 -745 -1891
rect -677 -1925 -665 -1891
rect -757 -1931 -665 -1925
rect -599 -1891 -507 -1885
rect -599 -1925 -587 -1891
rect -519 -1925 -507 -1891
rect -599 -1931 -507 -1925
rect -441 -1891 -349 -1885
rect -441 -1925 -429 -1891
rect -361 -1925 -349 -1891
rect -441 -1931 -349 -1925
rect -283 -1891 -191 -1885
rect -283 -1925 -271 -1891
rect -203 -1925 -191 -1891
rect -283 -1931 -191 -1925
rect -125 -1891 -33 -1885
rect -125 -1925 -113 -1891
rect -45 -1925 -33 -1891
rect -125 -1931 -33 -1925
rect 33 -1891 125 -1885
rect 33 -1925 45 -1891
rect 113 -1925 125 -1891
rect 33 -1931 125 -1925
rect 191 -1891 283 -1885
rect 191 -1925 203 -1891
rect 271 -1925 283 -1891
rect 191 -1931 283 -1925
rect 349 -1891 441 -1885
rect 349 -1925 361 -1891
rect 429 -1925 441 -1891
rect 349 -1931 441 -1925
rect 507 -1891 599 -1885
rect 507 -1925 519 -1891
rect 587 -1925 599 -1891
rect 507 -1931 599 -1925
rect 665 -1891 757 -1885
rect 665 -1925 677 -1891
rect 745 -1925 757 -1891
rect 665 -1931 757 -1925
rect 823 -1891 915 -1885
rect 823 -1925 835 -1891
rect 903 -1925 915 -1891
rect 823 -1931 915 -1925
rect 981 -1891 1073 -1885
rect 981 -1925 993 -1891
rect 1061 -1925 1073 -1891
rect 981 -1931 1073 -1925
rect 1139 -1891 1231 -1885
rect 1139 -1925 1151 -1891
rect 1219 -1925 1231 -1891
rect 1139 -1931 1231 -1925
rect -1287 -1975 -1241 -1963
rect -1287 -2351 -1281 -1975
rect -1247 -2351 -1241 -1975
rect -1287 -2363 -1241 -2351
rect -1129 -1975 -1083 -1963
rect -1129 -2351 -1123 -1975
rect -1089 -2351 -1083 -1975
rect -1129 -2363 -1083 -2351
rect -971 -1975 -925 -1963
rect -971 -2351 -965 -1975
rect -931 -2351 -925 -1975
rect -971 -2363 -925 -2351
rect -813 -1975 -767 -1963
rect -813 -2351 -807 -1975
rect -773 -2351 -767 -1975
rect -813 -2363 -767 -2351
rect -655 -1975 -609 -1963
rect -655 -2351 -649 -1975
rect -615 -2351 -609 -1975
rect -655 -2363 -609 -2351
rect -497 -1975 -451 -1963
rect -497 -2351 -491 -1975
rect -457 -2351 -451 -1975
rect -497 -2363 -451 -2351
rect -339 -1975 -293 -1963
rect -339 -2351 -333 -1975
rect -299 -2351 -293 -1975
rect -339 -2363 -293 -2351
rect -181 -1975 -135 -1963
rect -181 -2351 -175 -1975
rect -141 -2351 -135 -1975
rect -181 -2363 -135 -2351
rect -23 -1975 23 -1963
rect -23 -2351 -17 -1975
rect 17 -2351 23 -1975
rect -23 -2363 23 -2351
rect 135 -1975 181 -1963
rect 135 -2351 141 -1975
rect 175 -2351 181 -1975
rect 135 -2363 181 -2351
rect 293 -1975 339 -1963
rect 293 -2351 299 -1975
rect 333 -2351 339 -1975
rect 293 -2363 339 -2351
rect 451 -1975 497 -1963
rect 451 -2351 457 -1975
rect 491 -2351 497 -1975
rect 451 -2363 497 -2351
rect 609 -1975 655 -1963
rect 609 -2351 615 -1975
rect 649 -2351 655 -1975
rect 609 -2363 655 -2351
rect 767 -1975 813 -1963
rect 767 -2351 773 -1975
rect 807 -2351 813 -1975
rect 767 -2363 813 -2351
rect 925 -1975 971 -1963
rect 925 -2351 931 -1975
rect 965 -2351 971 -1975
rect 925 -2363 971 -2351
rect 1083 -1975 1129 -1963
rect 1083 -2351 1089 -1975
rect 1123 -2351 1129 -1975
rect 1083 -2363 1129 -2351
rect 1241 -1975 1287 -1963
rect 1241 -2351 1247 -1975
rect 1281 -2351 1287 -1975
rect 1241 -2363 1287 -2351
rect -1231 -2401 -1139 -2395
rect -1231 -2435 -1219 -2401
rect -1151 -2435 -1139 -2401
rect -1231 -2441 -1139 -2435
rect -1073 -2401 -981 -2395
rect -1073 -2435 -1061 -2401
rect -993 -2435 -981 -2401
rect -1073 -2441 -981 -2435
rect -915 -2401 -823 -2395
rect -915 -2435 -903 -2401
rect -835 -2435 -823 -2401
rect -915 -2441 -823 -2435
rect -757 -2401 -665 -2395
rect -757 -2435 -745 -2401
rect -677 -2435 -665 -2401
rect -757 -2441 -665 -2435
rect -599 -2401 -507 -2395
rect -599 -2435 -587 -2401
rect -519 -2435 -507 -2401
rect -599 -2441 -507 -2435
rect -441 -2401 -349 -2395
rect -441 -2435 -429 -2401
rect -361 -2435 -349 -2401
rect -441 -2441 -349 -2435
rect -283 -2401 -191 -2395
rect -283 -2435 -271 -2401
rect -203 -2435 -191 -2401
rect -283 -2441 -191 -2435
rect -125 -2401 -33 -2395
rect -125 -2435 -113 -2401
rect -45 -2435 -33 -2401
rect -125 -2441 -33 -2435
rect 33 -2401 125 -2395
rect 33 -2435 45 -2401
rect 113 -2435 125 -2401
rect 33 -2441 125 -2435
rect 191 -2401 283 -2395
rect 191 -2435 203 -2401
rect 271 -2435 283 -2401
rect 191 -2441 283 -2435
rect 349 -2401 441 -2395
rect 349 -2435 361 -2401
rect 429 -2435 441 -2401
rect 349 -2441 441 -2435
rect 507 -2401 599 -2395
rect 507 -2435 519 -2401
rect 587 -2435 599 -2401
rect 507 -2441 599 -2435
rect 665 -2401 757 -2395
rect 665 -2435 677 -2401
rect 745 -2435 757 -2401
rect 665 -2441 757 -2435
rect 823 -2401 915 -2395
rect 823 -2435 835 -2401
rect 903 -2435 915 -2401
rect 823 -2441 915 -2435
rect 981 -2401 1073 -2395
rect 981 -2435 993 -2401
rect 1061 -2435 1073 -2401
rect 981 -2441 1073 -2435
rect 1139 -2401 1231 -2395
rect 1139 -2435 1151 -2401
rect 1219 -2435 1231 -2401
rect 1139 -2441 1231 -2435
<< properties >>
string FIXED_BBOX -1378 -2520 1378 2520
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.5 m 8 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
