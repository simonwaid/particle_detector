magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< error_s >>
rect -331 -1140 -90 -1109
rect 230 -1140 471 -1109
rect -91 -1380 -90 -1349
rect 230 -1380 231 -1349
<< nwell >>
rect 1650 2620 1660 2790
<< pwell >>
rect -180 2030 850 2110
rect -1950 1380 -1780 1530
rect 670 1380 850 1530
rect -1950 860 -1750 920
rect 660 860 850 920
rect -1950 560 -1750 630
rect 660 560 850 620
rect -1950 -60 -1760 90
rect 690 -60 850 90
<< locali >>
rect -1910 3600 1710 3680
rect -190 2220 -80 3600
rect 1600 3050 1710 3600
rect 1600 2960 3780 3050
rect 1600 2220 1710 2400
rect 3530 2220 3780 2960
rect -2010 790 -1870 2130
rect 790 1260 920 2140
rect 1460 2110 3780 2220
rect 800 1010 920 1260
rect 1690 1800 3560 1890
rect 1690 1210 1790 1800
rect 3470 1230 3560 1800
rect 1670 1050 1780 1210
rect 790 790 920 1010
rect -2010 690 920 790
rect -2010 -640 -1870 690
rect 790 30 920 690
rect 1680 480 1780 1050
rect 3470 480 3560 1020
rect 1680 390 3560 480
rect 800 -640 910 30
rect -2010 -740 910 -640
rect -2010 -3330 -1870 -740
rect 720 -1180 910 -740
rect 720 -1360 730 -1180
rect 860 -1360 910 -1180
rect 720 -1500 910 -1360
rect 720 -1680 2700 -1500
<< viali >>
rect 1600 2400 1730 2960
rect 1590 1050 1670 1210
rect 3440 1020 3560 1230
rect 730 -1360 860 -1180
<< metal1 >>
rect -2000 3470 -1750 3540
rect -330 3470 60 3540
rect -2000 3000 -1850 3470
rect -180 3000 -100 3470
rect -2000 2830 1490 3000
rect 1594 2960 1736 2972
rect -2000 2360 -1850 2830
rect -180 2370 -100 2830
rect 1590 2400 1600 2960
rect 1730 2400 1740 2960
rect 1860 2830 3520 2870
rect 1594 2388 1736 2400
rect -2000 2290 -1750 2360
rect -330 2300 60 2370
rect 3480 2330 3520 2830
rect -2000 2070 -1850 2290
rect -180 2110 -100 2300
rect 1850 2290 3520 2330
rect -2000 2000 -1750 2070
rect -180 2030 930 2110
rect 660 2000 930 2030
rect -2000 1530 -1850 2000
rect 790 1530 930 2000
rect 1540 1550 1550 1740
rect 1800 1690 3340 1740
rect 1800 1680 1930 1690
rect 1800 1550 1820 1680
rect -2000 1380 930 1530
rect -2000 920 -1850 1380
rect 790 1210 930 1380
rect 1584 1210 1676 1222
rect 1730 1210 1820 1550
rect 3434 1230 3566 1242
rect 790 1050 840 1210
rect 1070 1050 1080 1210
rect 1580 1050 1590 1210
rect 1670 1050 1680 1210
rect 1730 1200 1910 1210
rect 1730 1080 3340 1200
rect 1730 1070 1910 1080
rect 790 920 930 1050
rect 1584 1038 1676 1050
rect -2000 860 -1750 920
rect 660 860 930 920
rect -2000 630 -1850 860
rect -2000 560 -1750 630
rect 790 620 930 860
rect 660 560 930 620
rect -2000 90 -1850 560
rect 790 90 930 560
rect 1730 600 1820 1070
rect 3430 1020 3440 1230
rect 3560 1020 3570 1230
rect 3434 1008 3566 1020
rect 1730 540 1910 600
rect -2000 -60 930 90
rect -2000 -530 -1850 -60
rect 790 -520 930 -60
rect 770 -530 930 -520
rect -2000 -580 -1750 -530
rect 660 -580 930 -530
rect -1960 -860 -1810 -800
rect -1960 -1330 -1860 -860
rect 724 -1180 866 -1168
rect -1960 -1480 -1810 -1330
rect 720 -1360 730 -1180
rect 860 -1360 870 -1180
rect 724 -1372 866 -1360
rect -1960 -1950 -1860 -1480
rect -1960 -2090 -1800 -1950
rect -1960 -2100 -1770 -2090
rect -1960 -2570 -1860 -2100
rect -1960 -2720 -1800 -2570
rect -1960 -3190 -1860 -2720
rect -1960 -3240 -1810 -3190
<< via1 >>
rect 1600 2400 1730 2960
rect 1550 1550 1800 1740
rect 840 1050 1070 1210
rect 1590 1050 1670 1210
rect 3440 1020 3560 1230
rect 730 -1360 860 -1180
<< metal2 >>
rect -1710 3420 1690 3440
rect -1710 3280 -260 3420
rect -20 3280 1690 3420
rect -1710 3270 1690 3280
rect 1440 3260 1690 3270
rect -1810 3190 1430 3200
rect -1810 3040 360 3190
rect 760 3040 1430 3190
rect -1810 3030 1430 3040
rect 1550 2980 1690 3260
rect 1550 2960 3280 2980
rect -1810 2790 1430 2800
rect -1810 2640 370 2790
rect 770 2640 1430 2790
rect -1810 2630 1430 2640
rect 1550 2570 1600 2960
rect 1440 2560 1600 2570
rect -1700 2540 1600 2560
rect -1700 2400 -260 2540
rect -20 2400 1600 2540
rect 1730 2620 3280 2960
rect 2220 2560 2660 2570
rect -300 2380 0 2400
rect 300 2390 340 2400
rect 1600 2390 1730 2400
rect 1800 2380 2220 2550
rect 2660 2380 3440 2550
rect 2220 2370 2660 2380
rect -90 1970 230 1980
rect -1710 1800 -90 1970
rect 230 1800 710 1970
rect -90 1790 230 1800
rect 1550 1740 1800 1750
rect -1800 1720 1550 1730
rect -1800 1570 370 1720
rect 770 1570 1550 1720
rect -1800 1560 1550 1570
rect 2220 1660 2660 1670
rect 1550 1540 1800 1550
rect 1850 1480 2220 1660
rect 2660 1480 3300 1660
rect 2220 1470 2660 1480
rect -1800 1350 770 1360
rect -1800 1200 370 1350
rect 1950 1240 3500 1420
rect -1800 1190 770 1200
rect 840 1210 1070 1220
rect 1590 1210 1670 1220
rect 1960 1210 2120 1240
rect 3310 1230 3560 1240
rect -190 1110 700 1120
rect -1710 360 -90 1110
rect 230 360 710 1110
rect 1070 1050 1590 1210
rect 1670 1050 2120 1210
rect 840 1040 1190 1050
rect 1590 1040 1670 1050
rect 1950 1040 2120 1050
rect 3390 1040 3440 1230
rect -180 350 310 360
rect -1810 280 770 290
rect -1810 130 370 280
rect -1810 120 770 130
rect -1800 -90 780 -80
rect -1800 -240 370 -90
rect 770 -240 780 -90
rect -1800 -250 780 -240
rect 980 -250 1190 1040
rect 1950 1020 3440 1040
rect 1950 1010 3560 1020
rect 1950 860 3500 1010
rect 2220 800 2660 810
rect 1850 620 2220 800
rect 2660 620 3300 800
rect 2220 610 2660 620
rect -90 -330 230 -320
rect -1710 -500 -90 -330
rect 230 -500 710 -330
rect -90 -510 230 -500
rect -760 -880 -440 -870
rect -1730 -1060 -760 -890
rect -440 -1060 770 -890
rect -760 -1070 -440 -1060
rect -1830 -1140 540 -1130
rect -1830 -1680 -90 -1140
rect 230 -1680 540 -1140
rect 630 -1170 770 -1060
rect 630 -1180 860 -1170
rect 630 -1360 730 -1180
rect 860 -1360 1050 -1180
rect 630 -1370 860 -1360
rect -90 -1690 230 -1680
rect 630 -1750 770 -1370
rect -1730 -1760 770 -1750
rect -1730 -2300 -760 -1760
rect -440 -2300 770 -1760
rect -760 -2310 -440 -2300
rect -1840 -2370 550 -2360
rect -1840 -2910 -90 -2370
rect 230 -2910 550 -2370
rect -90 -2920 230 -2910
rect -760 -2980 -440 -2970
rect 630 -2980 770 -2300
rect -1730 -3160 -760 -2980
rect -440 -3160 770 -2980
rect -760 -3170 -440 -3160
<< via2 >>
rect -260 3280 -20 3420
rect 360 3040 760 3190
rect 370 2640 770 2790
rect -260 2400 -20 2540
rect 2220 2380 2660 2560
rect -90 1800 230 1970
rect 370 1570 770 1720
rect 2220 1480 2660 1660
rect 370 1200 770 1350
rect -90 360 230 1110
rect 370 130 770 280
rect 370 -240 770 -90
rect 2220 620 2660 800
rect -90 -500 230 -330
rect -760 -1060 -440 -880
rect -90 -1680 230 -1140
rect -760 -2300 -440 -1760
rect -90 -2910 230 -2370
rect -760 -3160 -440 -2980
<< metal3 >>
rect -260 3430 -20 3440
rect -300 3090 -290 3430
rect 30 3090 40 3430
rect 360 3195 780 3200
rect 350 3190 780 3195
rect -260 2920 -20 3090
rect 350 3040 360 3190
rect 760 3040 780 3190
rect 350 3035 780 3040
rect -270 2760 -10 2920
rect 360 2790 780 3035
rect -260 2545 -20 2760
rect 360 2640 370 2790
rect 770 2640 780 2790
rect -270 2540 -10 2545
rect -270 2400 -260 2540
rect -20 2400 -10 2540
rect -270 2395 -10 2400
rect -100 1970 240 1975
rect -100 1800 -90 1970
rect 230 1800 240 1970
rect -100 1795 240 1800
rect -90 1115 230 1795
rect 360 1720 780 2640
rect 2210 2560 2670 2565
rect 2210 2380 2220 2560
rect 2660 2380 2670 2560
rect 2210 2375 2670 2380
rect 360 1570 370 1720
rect 770 1570 780 1720
rect 2220 1665 2660 2375
rect 360 1350 780 1570
rect 2210 1660 2670 1665
rect 2210 1480 2220 1660
rect 2660 1480 2670 1660
rect 2210 1475 2670 1480
rect 360 1200 370 1350
rect 770 1200 780 1350
rect 360 1195 780 1200
rect -100 1110 240 1115
rect -100 360 -90 1110
rect 230 360 240 1110
rect -100 355 240 360
rect 360 1010 770 1195
rect -90 -325 230 355
rect 360 280 780 1010
rect 2220 805 2660 1475
rect 2210 800 2670 805
rect 2210 620 2220 800
rect 2660 620 2670 800
rect 2210 615 2670 620
rect 360 130 370 280
rect 770 130 780 280
rect 360 -90 780 130
rect 360 -240 370 -90
rect 770 -240 780 -90
rect 360 -260 780 -240
rect -100 -330 240 -325
rect -100 -500 -90 -330
rect 230 -500 240 -330
rect -100 -505 240 -500
rect -770 -880 -430 -875
rect -770 -1060 -760 -880
rect -440 -1060 -430 -880
rect -770 -1065 -430 -1060
rect -760 -1220 -440 -1065
rect -90 -1135 230 -505
rect -100 -1140 240 -1135
rect -770 -1370 -430 -1220
rect -100 -1230 -90 -1140
rect -770 -1680 -760 -1370
rect -440 -1680 -430 -1370
rect -110 -1660 -90 -1230
rect -100 -1680 -90 -1660
rect 230 -1680 240 -1140
rect -760 -1755 -440 -1680
rect -100 -1685 240 -1680
rect -770 -1760 -430 -1755
rect -770 -2300 -760 -1760
rect -440 -2300 -430 -1760
rect -770 -2305 -430 -2300
rect -760 -2975 -440 -2305
rect -90 -2365 230 -1685
rect -100 -2370 240 -2365
rect -100 -2910 -90 -2370
rect 230 -2910 240 -2370
rect -100 -2915 240 -2910
rect -770 -2980 -430 -2975
rect -770 -3160 -760 -2980
rect -440 -3160 -430 -2980
rect -770 -3165 -430 -3160
<< via3 >>
rect -290 3420 30 3430
rect -290 3280 -260 3420
rect -260 3280 -20 3420
rect -20 3280 30 3420
rect -290 3090 30 3280
rect -760 -1680 -440 -1370
rect -90 -1670 230 -1350
<< metal4 >>
rect -291 3430 31 3431
rect -291 3090 -290 3430
rect 30 3090 31 3430
rect -291 3089 31 3090
rect -90 -1349 230 -960
rect -91 -1350 231 -1349
rect -761 -1370 -439 -1369
rect -761 -1680 -760 -1370
rect -440 -1680 -439 -1370
rect -91 -1670 -90 -1350
rect 230 -1670 231 -1350
rect -91 -1671 231 -1670
rect -761 -1681 -439 -1680
<< via4 >>
rect -290 3090 30 3430
rect -760 -1680 -440 -1370
<< metal5 >>
rect -320 3430 60 3460
rect -320 3090 -290 3430
rect 30 3090 60 3430
rect -320 2510 60 3090
rect -784 -1350 -416 -1346
rect -784 -1370 2950 -1350
rect -784 -1680 -760 -1370
rect -440 -1470 2950 -1370
rect -440 -1670 3760 -1470
rect -440 -1680 -416 -1670
rect -784 -1704 -416 -1680
rect 2610 -1790 3760 -1670
use dis_tran  dis_tran_0
timestamp 1654760956
transform 1 0 -1907 0 1 -3307
box -53 -53 2681 2621
use fb_transistor  fb_transistor_0
timestamp 1654760956
transform 1 0 -4020 0 1 -1780
box 5420 1880 7860 4782
use rf_transistors  rf_transistors_0
timestamp 1654760956
transform 1 0 -2380 0 1 2280
box 440 -2984 4042 1374
use sky130_fd_pr__cap_mim_m3_2_ZWVPUJ  sky130_fd_pr__cap_mim_m3_2_ZWVPUJ_0
timestamp 1654760956
transform 1 0 891 0 -1 760
box -2851 -1901 2873 1901
use tia_cur_mirror  tia_cur_mirror_0
timestamp 1654760956
transform 1 0 910 0 1 -660
box -60 -900 1822 740
<< end >>
