* SPICE3 file created from outd_stage3.ext - technology: sky130A

X0 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X15 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X16 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X39 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X40 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X41 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X42 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X43 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X45 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X48 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X51 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X53 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X56 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X57 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X58 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X59 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X61 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X64 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X65 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X66 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X67 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X69 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X70 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X72 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X75 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X76 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X77 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X80 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X83 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X85 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X90 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X92 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X93 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X94 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X98 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X99 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X100 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X101 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X102 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X104 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X105 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X106 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X107 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X108 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X109 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X110 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X111 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X112 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X113 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X114 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X115 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X116 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X117 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X118 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X119 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X120 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X121 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X122 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X123 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X124 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X125 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X126 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X127 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X128 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X129 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X130 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X131 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X132 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X133 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X134 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X135 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X136 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X137 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X138 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X139 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X140 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X141 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X142 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X143 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X145 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X146 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X147 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X148 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X149 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X150 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X151 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X152 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X153 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X154 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X155 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X156 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X157 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X158 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X159 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X160 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X161 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X162 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X163 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X164 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X165 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X166 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X167 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X168 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X169 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X170 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X171 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X172 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X173 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X174 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X175 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X176 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X177 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X178 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X179 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X180 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X181 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X182 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X183 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X184 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X185 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X186 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X187 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X188 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X189 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X190 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X191 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X192 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X193 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X194 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X195 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X196 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X197 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X198 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X199 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X200 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X201 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X202 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X203 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X204 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X205 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X206 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X207 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X208 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X209 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X210 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X211 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X212 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X213 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X214 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X215 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X216 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X217 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X218 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X219 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X220 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X221 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X222 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X223 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X224 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X225 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X226 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X227 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X228 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X229 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X230 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X231 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X232 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X233 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X234 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X235 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X236 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X237 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X238 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X239 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X240 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X241 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X242 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X243 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X244 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X245 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X246 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X247 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X248 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X249 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X250 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X251 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X252 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X253 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X254 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X255 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X256 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X257 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X258 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X259 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X261 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X262 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X263 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X264 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X265 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X266 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X267 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X268 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X269 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X273 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X274 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X275 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X276 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X277 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X279 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X280 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X281 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X283 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X284 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X285 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X286 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X287 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X288 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X289 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X290 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X291 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X292 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X293 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X294 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X295 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X296 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X297 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X298 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X299 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X300 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X301 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X302 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X303 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X304 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X305 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X306 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X307 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X308 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X309 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X310 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X311 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X312 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X313 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X314 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X315 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X316 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X317 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X318 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X319 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X320 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X321 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X322 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X323 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X324 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X325 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X326 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X327 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X328 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X329 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X330 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X331 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X332 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X333 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X334 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X335 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X336 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X337 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X338 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X339 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X340 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X341 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X342 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X343 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X344 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X345 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X346 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X347 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X348 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X349 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X350 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X351 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X352 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X353 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X354 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X355 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X356 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X357 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X358 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X359 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X360 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X361 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X362 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X363 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X364 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X365 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X366 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X367 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X368 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X369 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X370 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X371 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X372 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X373 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X374 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X375 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X376 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X377 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X378 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X379 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X380 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X381 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X382 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X383 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X384 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X385 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X386 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X387 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X388 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X389 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X390 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X391 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X392 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X393 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X394 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X395 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X396 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X397 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X398 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X399 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X400 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X401 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X402 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X403 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X404 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X405 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X406 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X407 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X408 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X409 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X410 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X411 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X412 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X413 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X414 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X415 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X416 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X417 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X418 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X419 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X420 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X421 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X422 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X423 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X424 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X425 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X426 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X427 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X428 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X429 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X430 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X431 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X432 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X433 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X434 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X435 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X436 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X437 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X438 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X439 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X440 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X441 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X442 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X443 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X444 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X445 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X446 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X447 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X448 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X449 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X450 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X451 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X452 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X453 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X454 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X455 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X456 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X457 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X458 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X459 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X460 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X461 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X462 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X463 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X464 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X465 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X466 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X467 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X468 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X469 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X470 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X471 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X472 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X473 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X474 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X475 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X476 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X477 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X478 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X479 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X480 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X481 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X482 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X483 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X484 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X485 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X486 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X487 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X488 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X489 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X490 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X491 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X492 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X493 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X494 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X495 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X496 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X497 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X498 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X499 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X500 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X501 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X502 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X503 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X504 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X505 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X506 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X507 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X508 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X509 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X510 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X511 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X512 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X513 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X514 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X515 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X516 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X517 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X519 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X520 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X521 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X522 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X523 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X524 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X525 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X526 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X527 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X528 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X529 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X530 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X531 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X532 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X533 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X534 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X535 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X536 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X537 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X538 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X540 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X541 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X542 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X543 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X544 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X545 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X546 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X547 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X548 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X549 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X550 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X551 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X552 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X553 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X554 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X555 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X556 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X557 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X558 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X559 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X560 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X561 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X562 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X563 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X564 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X565 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X566 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X567 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X568 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X569 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X570 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X571 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X572 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X573 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X574 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X575 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X576 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X577 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X578 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X579 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X580 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X581 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X582 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X583 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X584 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X585 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X586 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X587 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X588 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X589 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X590 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X591 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X592 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X593 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X594 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X595 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X596 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X597 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X598 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X599 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X600 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X601 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X602 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X603 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X604 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X605 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X606 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X607 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X608 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X609 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X610 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X611 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X612 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X613 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X614 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X615 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X616 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X617 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X618 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X619 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X620 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X621 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X622 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X623 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X624 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X625 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X626 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X627 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X628 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X629 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X630 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X631 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X632 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X633 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X634 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X635 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X636 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X637 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X638 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X639 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X640 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X641 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X642 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X643 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X644 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X645 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X646 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X647 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X648 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X649 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X650 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X651 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X652 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X653 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X654 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X655 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X656 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X657 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X658 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X659 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X660 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X661 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X662 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X663 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X664 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X665 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X666 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X667 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X668 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X669 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X670 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X671 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X672 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X673 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X674 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X675 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X676 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X677 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X678 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X679 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X680 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X681 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X682 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X683 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X684 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X685 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X686 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X687 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X688 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X689 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X690 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X691 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X692 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X693 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X694 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X695 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X696 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X697 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X698 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X699 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X700 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X701 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X702 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X703 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X704 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X705 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X706 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X707 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X708 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X709 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X710 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X711 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X712 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X713 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X714 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X715 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X716 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X717 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X718 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X719 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X720 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X721 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X722 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X723 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X724 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X725 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X726 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X727 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X728 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X729 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X730 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X731 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X732 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X733 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X734 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X735 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X736 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X737 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X738 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X739 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X740 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X741 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X742 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X743 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X744 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X745 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X746 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X747 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X748 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X749 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X750 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X751 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X752 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X753 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X754 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X755 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X756 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X757 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X758 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X759 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X760 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X761 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X762 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X763 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X764 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X765 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X766 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X767 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X768 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X769 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X770 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X771 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X772 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X773 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X774 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X775 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X776 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X777 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X778 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X779 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X780 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X781 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X782 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X783 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X784 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X785 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X786 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X787 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X788 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X789 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X790 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X791 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X792 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X793 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X794 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X795 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X796 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X797 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X798 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X799 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X800 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X801 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X802 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X803 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X804 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X805 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X806 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X807 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X808 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X809 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X810 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X811 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X812 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X813 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X814 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X815 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X816 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X817 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X818 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X819 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X820 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X821 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X822 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X823 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X824 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X825 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X826 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X827 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X828 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X829 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X830 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X831 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X832 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X833 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X834 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X835 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X836 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X837 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X838 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X839 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X840 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X841 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X842 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X843 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X844 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X845 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X846 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X847 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X848 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X849 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X850 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X851 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X852 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X853 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X854 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X855 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X856 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X857 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X858 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X859 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X860 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X861 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X862 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X863 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X864 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X865 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X866 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X867 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X868 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X869 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X870 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X871 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X872 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X873 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X874 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X875 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X876 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X877 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X878 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X879 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X880 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X881 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X882 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X883 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X884 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X885 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X886 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X887 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X888 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X889 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X890 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X891 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X892 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X893 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X894 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X895 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X896 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X897 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X898 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X899 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X900 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X901 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X902 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X903 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X904 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X905 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X906 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X907 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X908 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X909 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X910 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X911 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X912 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X913 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X914 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X915 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X916 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X917 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X918 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X919 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X920 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X921 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X922 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X923 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X924 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X925 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X926 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X927 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X928 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X929 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X930 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X931 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X932 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X933 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X934 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X935 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X936 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X937 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X938 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X939 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X940 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X941 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X942 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X943 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X944 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X945 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X946 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X947 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X948 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X949 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X950 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X951 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X952 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X953 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X954 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X955 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X956 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X957 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X958 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X959 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X960 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X961 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X962 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X963 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X964 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X965 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X966 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X967 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X968 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X969 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X970 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X971 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X972 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X973 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X974 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X975 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X976 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X977 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X978 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X979 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X980 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X981 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X982 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X983 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X984 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X985 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X986 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X987 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X988 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X989 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X990 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X991 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X992 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X993 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X994 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X995 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X996 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X997 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X998 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X999 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1000 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1001 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1002 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1003 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1004 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1005 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1006 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1007 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1008 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1009 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1010 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1011 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1012 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1013 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1014 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1015 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1016 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1017 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1018 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1019 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1020 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1021 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1022 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1023 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1024 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1025 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1026 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1027 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1028 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1029 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1030 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1031 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1032 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1033 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1034 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1035 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1036 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1037 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1038 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1039 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1040 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1041 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1042 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1043 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1044 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1045 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1046 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1047 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1048 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1049 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1050 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1051 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1052 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1053 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1054 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1055 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1056 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1057 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1058 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1059 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1060 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1061 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1062 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1063 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1064 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1065 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1066 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1067 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1068 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1069 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1070 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1071 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1072 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1073 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1074 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1075 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1076 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1077 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1078 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1079 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1080 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1081 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1082 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1083 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1084 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1085 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1086 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1087 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1088 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1089 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1090 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1091 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1092 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1093 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1094 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1095 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1096 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1097 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1098 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1099 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1100 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1101 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1102 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1103 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1104 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1105 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1106 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1107 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1108 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1109 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1110 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1111 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1112 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1113 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1114 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1115 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1116 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1117 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1118 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1119 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1120 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1121 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1122 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1123 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1124 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1125 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1126 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1127 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1128 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1129 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1130 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1131 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1132 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1133 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1134 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1135 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1136 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1137 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1138 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1139 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1140 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1141 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1142 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1143 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1144 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1145 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1146 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1147 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1148 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1149 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1150 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1151 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1152 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1153 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1154 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1155 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1156 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1157 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1158 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1159 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1160 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1161 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1162 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1163 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1164 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1165 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1166 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1167 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1168 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1169 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1170 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1171 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1172 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1173 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1174 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1175 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1176 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1177 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1178 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1179 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1180 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1181 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1182 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1183 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1184 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1185 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1186 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1187 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1188 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1189 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1190 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1191 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1192 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1193 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1194 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1195 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1196 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1197 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1198 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1199 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1200 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1201 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1202 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1203 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1204 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1205 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1206 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1207 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1208 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1209 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1210 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1211 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1212 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1213 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1214 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1215 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1216 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1217 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1218 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1219 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1220 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1221 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1222 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1223 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1224 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1225 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1226 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1227 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1228 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1229 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1230 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1231 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1232 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1233 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1234 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1235 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1236 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1237 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1238 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1239 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1240 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1241 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1242 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1243 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1244 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1245 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1246 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1247 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1248 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1249 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1250 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1251 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1252 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1253 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1254 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1255 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1256 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1257 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1258 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1259 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1260 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1261 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1262 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1263 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1264 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1265 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1266 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1267 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1268 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1269 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1270 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1271 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1272 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1273 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1274 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1275 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1276 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1277 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1278 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1279 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1280 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1281 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1282 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1283 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1284 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1285 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1286 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1287 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1288 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1289 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1290 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1291 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1292 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1293 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1294 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1295 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1296 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1297 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1298 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1299 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1300 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1301 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1302 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1303 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1304 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1305 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1306 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1307 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1308 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1309 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1310 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1311 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1312 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1313 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1314 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1315 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1316 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1317 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1318 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1319 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1320 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1321 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1322 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1323 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1324 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1325 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1326 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1327 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1328 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1329 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1330 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1331 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1332 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1333 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1334 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1335 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1336 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1337 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1338 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1339 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1340 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1341 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1342 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1343 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1344 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1345 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1346 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1347 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1348 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1349 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1350 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1351 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1352 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1353 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1354 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1355 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1356 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1357 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1358 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1359 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1360 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1361 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1362 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1363 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1364 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1365 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1366 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1367 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1368 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1369 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1370 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1371 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1372 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1373 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1374 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1375 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1376 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1377 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1378 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1379 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1380 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1381 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1382 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1383 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1384 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1385 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1386 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1387 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1388 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1389 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1390 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1391 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1392 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1393 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1394 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1395 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1396 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1397 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1398 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1399 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1400 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1401 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1402 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1403 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1404 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1405 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1406 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1407 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1408 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1409 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1410 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1411 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1412 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1413 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1414 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1415 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1416 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1417 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1418 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1419 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1420 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1421 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1422 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1423 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1424 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1425 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1426 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1427 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1428 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1429 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1430 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1431 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1432 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1433 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1434 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1435 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1436 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1437 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1438 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1439 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1440 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1441 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1442 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1443 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1444 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1445 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1446 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1447 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1448 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1449 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1450 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1451 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1452 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1453 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1454 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1455 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1456 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1457 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1458 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1459 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1460 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1461 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1462 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1463 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1464 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1465 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1466 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1467 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1468 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1469 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1470 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1471 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1472 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1473 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1474 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1475 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1476 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1477 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1478 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1479 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1480 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1481 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1482 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1483 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1484 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1485 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1486 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1487 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1488 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1489 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1490 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1491 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1492 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1493 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1494 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1495 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1496 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1497 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1498 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1499 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1500 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1501 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1502 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1503 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1504 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1505 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1506 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1507 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1508 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1509 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1510 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1511 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1512 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1513 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1514 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1515 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1516 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1517 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1518 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1519 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1520 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1521 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1522 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1523 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1524 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1525 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1526 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1527 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1528 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1529 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1530 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1531 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1532 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1533 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1534 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1535 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1536 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1537 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1538 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1539 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1540 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1541 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1542 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1543 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1544 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1545 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1546 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1547 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1548 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1549 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1550 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1551 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1552 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1553 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1554 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1555 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1556 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1557 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1558 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1559 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1560 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1561 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1562 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1563 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1564 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1565 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1566 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1567 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1568 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1569 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1570 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1571 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1572 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1573 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1574 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1575 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1576 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1577 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1578 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1579 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1580 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1581 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1582 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1583 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1584 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1585 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1586 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1587 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1588 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1589 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1590 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1591 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1592 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1593 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1594 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1595 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1596 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1597 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1598 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1599 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1600 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1601 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1602 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1603 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1604 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1605 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1606 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1607 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1608 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1609 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1610 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1611 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1612 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1613 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1614 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1615 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1616 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1617 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1618 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1619 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1620 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1621 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1622 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1623 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1624 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1625 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1626 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1627 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1628 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1629 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1630 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1631 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1632 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1633 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1634 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1635 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1636 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1637 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1638 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1639 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1640 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1641 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1642 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1643 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1644 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1645 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1646 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1647 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1648 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1649 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1650 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1651 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1652 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1653 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1654 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1655 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1656 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1657 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1658 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1659 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1660 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1661 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1662 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1663 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1664 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1665 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1666 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1667 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1668 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1669 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1670 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1671 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1672 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1673 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1674 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1675 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1676 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1677 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1678 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1679 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1680 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1681 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1682 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1683 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1684 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1685 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1686 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1687 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1688 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1689 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1690 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1691 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1692 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1693 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1694 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1695 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1696 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1697 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1698 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1699 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1700 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1701 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1702 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1703 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1704 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1705 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1706 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1707 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1708 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1709 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1710 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1711 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1712 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1713 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1714 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1715 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1716 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1717 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1718 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1719 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1720 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1721 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1722 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1723 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1724 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1725 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1726 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1727 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1728 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1729 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1730 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1731 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1732 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1733 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1734 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1735 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1736 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1737 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1738 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1739 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1740 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1741 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1742 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1743 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1744 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1745 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1746 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1747 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1748 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1749 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1750 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1751 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1752 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1753 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1754 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1755 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1756 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1757 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1758 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1759 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1760 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1761 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1762 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1763 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1764 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1765 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1766 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1767 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1768 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1769 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1770 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1771 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1772 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1773 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1774 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1775 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1776 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1777 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1778 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1779 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1780 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1781 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1782 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1783 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1784 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1785 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1786 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1787 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1788 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1789 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1790 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1791 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1792 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1793 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1794 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1795 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1796 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1797 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1798 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1799 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1800 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1801 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1802 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1803 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1804 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1805 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1806 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1807 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1808 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1809 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1810 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1811 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1812 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1813 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1814 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1815 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1816 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1817 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1818 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1819 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1820 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1821 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1822 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1823 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1824 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1825 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1826 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1827 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1828 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1829 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1830 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1831 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1832 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1833 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1834 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1835 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1836 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1837 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1838 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1839 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1840 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1841 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1842 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1843 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1844 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1845 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1846 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1847 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1848 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1849 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1850 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1851 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1852 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1853 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1854 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1855 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1856 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1857 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1858 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1859 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1860 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1861 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1862 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1863 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1864 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1865 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1866 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1867 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1868 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1869 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1870 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1871 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1872 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1873 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1874 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1875 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1876 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1877 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1878 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1879 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1880 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1881 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1882 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1883 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1884 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1885 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1886 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1887 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1888 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1889 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1890 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1891 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1892 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1893 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1894 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1895 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1896 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1897 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1898 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1899 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1900 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1901 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1902 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1903 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1904 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1905 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1906 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1907 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1908 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1909 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1910 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1911 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1912 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1913 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1914 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1915 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1916 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1917 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1918 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1919 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1920 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1921 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1922 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1923 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1924 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1925 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1926 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1927 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1928 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1929 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1930 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1931 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1932 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1933 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1934 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1935 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1936 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1937 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1938 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1939 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1940 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1941 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1942 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1943 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1944 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1945 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1946 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1947 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1948 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1949 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1950 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1951 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1952 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1953 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1954 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1955 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1956 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1957 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1958 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1959 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1960 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1961 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1962 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1963 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1964 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1965 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1966 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1967 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1968 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1969 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1970 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1971 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1972 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1973 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1974 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1975 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1976 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1977 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1978 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1979 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1980 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1981 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1982 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1983 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1984 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1985 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1986 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1987 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1988 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1989 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1990 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1991 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1992 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1993 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1994 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1995 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1996 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1997 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1998 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1999 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2000 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2001 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2002 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2003 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2004 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2005 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2006 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2007 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2008 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2009 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2010 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2011 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2012 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2013 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2014 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2015 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2016 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2017 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2018 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2019 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2020 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2021 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2022 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2023 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2024 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2025 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2026 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2027 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2028 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2029 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2030 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2031 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2032 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2033 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2034 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2035 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2036 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2037 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2038 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2039 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2040 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2041 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2042 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2043 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2044 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2045 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2046 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2047 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2048 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2049 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2050 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2051 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2052 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2053 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2054 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2055 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2056 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2057 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2058 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2059 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2060 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2061 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2062 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2063 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2064 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2065 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2066 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2067 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2068 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2069 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2070 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2071 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2072 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2073 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2074 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2075 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2076 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2077 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2078 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2079 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2080 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2081 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2082 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2083 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2084 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2085 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2086 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2087 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2088 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2089 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2090 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2091 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2092 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2093 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2094 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2095 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2096 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2097 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2098 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2099 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2100 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2101 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2102 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2103 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2104 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2105 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2106 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2107 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2108 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2109 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2110 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2111 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2112 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2113 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2114 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2115 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2116 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2117 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2118 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2119 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2120 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2121 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2122 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2123 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2124 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2125 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2126 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2127 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2128 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2129 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2130 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2131 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2132 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2133 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2134 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2135 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2136 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2137 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2138 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2139 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2140 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2141 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2142 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2143 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2144 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2145 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2146 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2147 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2148 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2149 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2150 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2151 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2152 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2153 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2154 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2155 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2156 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2157 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2158 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2159 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2160 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2161 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2162 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2163 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2164 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2165 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2166 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2167 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2168 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2169 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2170 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2171 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2172 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2173 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2174 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2175 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2176 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2177 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2178 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2179 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2180 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2181 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2182 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2183 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2184 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2185 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2186 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2187 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2188 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2189 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2190 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2191 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2192 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2193 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2194 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2195 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2196 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2197 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2198 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2199 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2200 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2201 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2202 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2203 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2204 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2205 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2206 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2207 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2208 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2209 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2210 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2211 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2212 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2213 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2214 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2215 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2216 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2217 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2218 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2219 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2220 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2221 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2222 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2223 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2224 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2225 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2226 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2227 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2228 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2229 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2230 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2231 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2232 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2233 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2234 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2235 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2236 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2237 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2238 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2239 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2240 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2241 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2242 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2243 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2244 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2245 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2246 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2247 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2248 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2249 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2250 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2251 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2252 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2253 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2254 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2255 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2256 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2257 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2258 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2259 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2260 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2261 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2262 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2263 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2264 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2265 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2266 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2267 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2268 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2269 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2270 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2271 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2272 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2273 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2274 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2275 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2276 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2277 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2278 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2279 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2280 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2281 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2282 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2283 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2284 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2285 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2286 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2287 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2288 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2289 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2290 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2291 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2292 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2293 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2294 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2295 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2296 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2297 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2298 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2299 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2300 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2301 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2302 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2303 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2304 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2305 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2306 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2307 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2308 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2309 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2310 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2311 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2312 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2313 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2314 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2315 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2316 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2317 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2318 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2319 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2320 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2321 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2322 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2323 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2324 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2325 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2326 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2327 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2328 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2329 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2330 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2331 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2332 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2333 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2334 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2335 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2336 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2337 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2338 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2339 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2340 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2341 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2342 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2343 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2344 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2345 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2346 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2347 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2348 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2349 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2350 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2351 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2352 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2353 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2354 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2355 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2356 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2357 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2358 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2359 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2360 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2361 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2362 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2363 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2364 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2365 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2366 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2367 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2368 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2369 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2370 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2371 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2372 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2373 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2374 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2375 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2376 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2377 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2378 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2379 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2380 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2381 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2382 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2383 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2384 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2385 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2386 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2387 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2388 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2389 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2390 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2391 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2392 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2393 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2394 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2395 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2396 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2397 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2398 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2399 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2400 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2401 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2402 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2403 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2404 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2405 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2406 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2407 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2408 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2409 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2410 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2411 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2412 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2413 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2414 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2415 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2416 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2417 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2418 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2419 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2420 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2421 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2422 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2423 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2424 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2425 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2426 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2427 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2428 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2429 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2430 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2431 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2432 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2433 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2434 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2435 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2436 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2437 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2438 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2439 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2440 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2441 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2442 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2443 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2444 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2445 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2446 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2447 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2448 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2449 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2450 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2451 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2452 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2453 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2454 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2455 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2456 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2457 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2458 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2459 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2460 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2461 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2462 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2463 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2464 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2465 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2466 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2467 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2468 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2469 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2470 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2471 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2472 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2473 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2474 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2475 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2476 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2477 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2478 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2479 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2480 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2481 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2482 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2483 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2484 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2485 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2486 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2487 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2488 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2489 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2490 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2491 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2492 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2493 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2494 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2495 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2496 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2497 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2498 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2499 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2500 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2501 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2502 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2503 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2504 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2505 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2506 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2507 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2508 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2509 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2510 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2511 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2512 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2513 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2514 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2515 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2516 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2517 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2518 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2519 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2520 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2521 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2522 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2523 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2524 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2525 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2526 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2527 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2528 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2529 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2530 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2531 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2532 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2533 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2534 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2535 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2536 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2537 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2538 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2539 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2540 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2541 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2542 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2543 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2544 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2545 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2546 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2547 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2548 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2549 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2550 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2551 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2552 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2553 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2554 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2555 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2556 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2557 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2558 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2559 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2560 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2561 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2562 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2563 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2564 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2565 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2566 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2567 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2568 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2569 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2570 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2571 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2572 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2573 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2574 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2575 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2576 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2577 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2578 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2579 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2580 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2581 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2582 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2583 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2584 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2585 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2586 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2587 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2588 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2589 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2590 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2591 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2592 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2593 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2594 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2595 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2596 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2597 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2598 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2599 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2600 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2601 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2602 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2603 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2604 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2605 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2606 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2607 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2608 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2609 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2610 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2611 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2612 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2613 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2614 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2615 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2616 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2617 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2618 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2619 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2620 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2621 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2622 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2623 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2624 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2625 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2626 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2627 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2628 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2629 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2630 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2631 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2632 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2633 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2634 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2635 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2636 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2637 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2638 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2639 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2640 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2641 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2642 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2643 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2644 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2645 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2646 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2647 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2648 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2649 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2650 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2651 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2652 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2653 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2654 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2655 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2656 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2657 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2658 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2659 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2660 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2661 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2662 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2663 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2664 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2665 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2666 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2667 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2668 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2669 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2670 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2671 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2672 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2673 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2674 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2675 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2676 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2677 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2678 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2679 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2680 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2681 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2682 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2683 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2684 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2685 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2686 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2687 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2688 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2689 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2690 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2691 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2692 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2693 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2694 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2695 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2696 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2697 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2698 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2699 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2700 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2701 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2702 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2703 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2704 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2705 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2706 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2707 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2708 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2709 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2710 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2711 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2712 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2713 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2714 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2715 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2716 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2717 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2718 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2719 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2720 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2721 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2722 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2723 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2724 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2725 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2726 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2727 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2728 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2729 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2730 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2731 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2732 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2733 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2734 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2735 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2736 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2737 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2738 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2739 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2740 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2741 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2742 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2743 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2744 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2745 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2746 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2747 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2748 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2749 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2750 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2751 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2752 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2753 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2754 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2755 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2756 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2757 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2758 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2759 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2760 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2761 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2762 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2763 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2764 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2765 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2766 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2767 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2768 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2769 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2770 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2771 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2772 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2773 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2774 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2775 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2776 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2777 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2778 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2779 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2780 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2781 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2782 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2783 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2784 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2785 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2786 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2787 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2788 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2789 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2790 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2791 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2792 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2793 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2794 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2795 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2796 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2797 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2798 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2799 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2800 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2801 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2802 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2803 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2804 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2805 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2806 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2807 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2808 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2809 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2810 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2811 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2812 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2813 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2814 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2815 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2816 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2817 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2818 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2819 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2820 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2821 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2822 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2823 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2824 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2825 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2826 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2827 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2828 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2829 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2830 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2831 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2832 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2833 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2834 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2835 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2836 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2837 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2838 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2839 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2840 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2841 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2842 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2843 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2844 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2845 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2846 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2847 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2848 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2849 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2850 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2851 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2852 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2853 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2854 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2855 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2856 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2857 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2858 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2859 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2860 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2861 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2862 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2863 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2864 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2865 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2866 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2867 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2868 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2869 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2870 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2871 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2872 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2873 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2874 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2875 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2876 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2877 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2878 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2879 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2880 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2881 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2882 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2883 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2884 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2885 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2886 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2887 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2888 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2889 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2890 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2891 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2892 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2893 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2894 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2895 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2896 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2897 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2898 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2899 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2900 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2901 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2902 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2903 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2904 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2905 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2906 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2907 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2908 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2909 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2910 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2911 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2912 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2913 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2914 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2915 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2916 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2917 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2918 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2919 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2920 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2921 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2922 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2923 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2924 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2925 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2926 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2927 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2928 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2929 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2930 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2931 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2932 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2933 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2934 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2935 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2936 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2937 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2938 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2939 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2940 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2941 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2942 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2943 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2944 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2945 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2946 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2947 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2948 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2949 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2950 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2951 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2952 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2953 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2954 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2955 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2956 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2957 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2958 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2959 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2960 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2961 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2962 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2963 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2964 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2965 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2966 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2967 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2968 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2969 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2970 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2971 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2972 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2973 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2974 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2975 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2976 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2977 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2978 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2979 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2980 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2981 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2982 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2983 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2984 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2985 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2986 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2987 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2988 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2989 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2990 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2991 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2992 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2993 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2994 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2995 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2996 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2997 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2998 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2999 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3000 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3001 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3002 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3003 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3004 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3005 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3006 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3007 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3008 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3009 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3010 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3011 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3012 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3013 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3014 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3015 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3016 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3017 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3018 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3019 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3020 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3021 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3022 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3023 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3024 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3025 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3026 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3027 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3028 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3029 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3030 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3031 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3032 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3033 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3034 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3035 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3036 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3037 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3038 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3039 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3040 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3041 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3042 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3043 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3044 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3045 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3046 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3047 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3048 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3049 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3050 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3051 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3052 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3053 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3054 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3055 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3056 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3057 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3058 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3059 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3060 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3061 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3062 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3063 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3064 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3065 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3066 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3067 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3068 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3069 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3070 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3071 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3072 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3073 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3074 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3075 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3076 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3077 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3078 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3079 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3080 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3081 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3082 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3083 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3084 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3085 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3086 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3087 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3088 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3089 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3090 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3091 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3092 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3093 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3094 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3095 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3096 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3097 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3098 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3099 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3100 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3101 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3102 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3103 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3104 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3105 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3106 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3107 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3108 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3109 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3110 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3111 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3112 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3113 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3114 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3115 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3116 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3117 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3118 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3119 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3120 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3121 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3122 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3123 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3124 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3125 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3126 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3127 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3128 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3129 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3130 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3131 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3132 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3133 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3134 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3135 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3136 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3137 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3138 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3139 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3140 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3141 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3142 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3143 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3144 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3145 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3146 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3147 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3148 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3149 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3150 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3151 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3152 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3153 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3154 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3155 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3156 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3157 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3158 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3159 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3160 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3161 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3162 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3163 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3164 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3165 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3166 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3167 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3168 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3169 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3170 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3171 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3172 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3173 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3174 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3175 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3176 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3177 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3178 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3179 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3180 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3181 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3182 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3183 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3184 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3185 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3186 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3187 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3188 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3189 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3190 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3191 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3192 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3193 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3194 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3195 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3196 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3197 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3198 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3199 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3200 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3201 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3202 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3203 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3204 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3205 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3206 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3207 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3208 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3209 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3210 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3211 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3212 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3213 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3214 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3215 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3216 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3217 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3218 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3219 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3220 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3221 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3222 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3223 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3224 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3225 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3226 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3227 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3228 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3229 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3230 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3231 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3232 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3233 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3234 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3235 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3236 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3237 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3238 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3239 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3240 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3241 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3242 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3243 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3244 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3245 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3246 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3247 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3248 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3249 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3250 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3251 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3252 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3253 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3254 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3255 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3256 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3257 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3258 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3259 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3260 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3261 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3262 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3263 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3264 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3265 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3266 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3267 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3268 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3269 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3270 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3271 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3272 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3273 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3274 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3275 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3276 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3277 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3278 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3279 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3280 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3281 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3282 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3283 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3284 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3285 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3286 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3287 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3288 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3289 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3290 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3291 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3292 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3293 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3294 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3295 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3296 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3297 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3298 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3299 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3300 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3301 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3302 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3303 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3304 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3305 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3306 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3307 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3308 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3309 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3310 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3311 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3312 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3313 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3314 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3315 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3316 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3317 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3318 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3319 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3320 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3321 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3322 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3323 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3324 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3325 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3326 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3327 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3328 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3329 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3330 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3331 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3332 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3333 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3334 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3335 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3336 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3337 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3338 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3339 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3340 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3341 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3342 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3343 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3344 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3345 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3346 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3347 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3348 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3349 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3350 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3351 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3352 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3353 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3354 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3355 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3356 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3357 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3358 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3359 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3360 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3361 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3362 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3363 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3364 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3365 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3366 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3367 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3368 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3369 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3370 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3371 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3372 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3373 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3374 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3375 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3376 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3377 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3378 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3379 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3380 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3381 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3382 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3383 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3384 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3385 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3386 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3387 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3388 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3389 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3390 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3391 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3392 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3393 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3394 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3395 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3396 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3397 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3398 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3399 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3400 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3401 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3402 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3403 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3404 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3405 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3406 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3407 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3408 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3409 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3410 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3411 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3412 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3413 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3414 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3415 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3416 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3417 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3418 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3419 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3420 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3421 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3422 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3423 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3424 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3425 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3426 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3427 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3428 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3429 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3430 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3431 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3432 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3433 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3434 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3435 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3436 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3437 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3438 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3439 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3440 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3441 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3442 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3443 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3444 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3445 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3446 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3447 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3448 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3449 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3450 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3451 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3452 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3453 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3454 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3455 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3456 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3457 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3458 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3459 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3460 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3461 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3462 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3463 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3464 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3465 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3466 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3467 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3468 m3_11690_14240# m4_40470_12200# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3469 m3_11690_14240# m4_40470_12880# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3470 m4_40470_12880# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3471 m4_40470_12200# m3_11690_14240# VSUBS sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3472 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3473 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3474 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3475 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3476 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3477 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3478 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3479 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3480 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3481 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3482 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3483 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3484 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3485 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3486 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3487 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3488 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3489 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3490 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3491 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3492 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3493 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3494 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3495 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3496 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3497 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3498 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3499 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3500 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3501 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3502 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3503 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3504 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3505 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3506 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3507 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3508 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3509 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3510 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3511 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3512 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3513 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3514 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3515 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3516 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3517 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3518 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3519 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3520 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3521 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3522 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3523 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3524 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3525 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3526 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3527 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3528 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3529 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3530 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3531 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3532 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3533 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3534 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3535 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3536 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3537 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3538 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3539 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3540 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3541 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3542 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3543 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3544 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3545 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3546 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3547 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3548 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3549 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3550 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3551 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3552 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3553 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3554 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3555 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3556 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3557 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3558 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3559 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3560 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3561 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3562 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3563 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3564 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3565 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3566 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3567 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3568 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3569 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3570 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3571 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3572 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3573 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3574 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3575 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3576 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3577 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3578 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3579 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3580 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3581 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3582 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3583 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3584 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3585 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3586 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3587 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3588 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3589 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3590 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3591 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3592 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3593 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3594 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3595 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3596 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3597 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3598 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3599 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3600 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3601 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3602 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3603 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3604 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3605 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3606 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3607 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3608 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3609 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3610 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3611 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3612 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3613 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3614 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3615 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3616 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3617 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3618 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3619 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3620 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3621 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3622 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3623 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3624 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3625 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3626 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3627 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3628 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3629 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3630 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3631 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3632 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3633 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3634 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3635 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3636 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3637 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3638 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3639 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3640 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3641 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3642 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3643 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3644 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3645 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3646 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3647 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3648 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3649 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3650 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3651 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3652 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3653 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3654 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3655 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3656 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3657 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3658 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3659 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3660 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3661 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3662 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3663 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3664 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3665 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3666 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3667 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3668 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3669 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3670 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3671 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3672 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3673 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3674 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3675 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3676 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3677 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3678 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3679 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3680 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3681 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3682 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3683 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3684 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3685 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3686 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3687 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3688 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3689 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3690 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3691 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3692 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3693 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3694 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3695 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3696 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3697 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3698 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3699 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3700 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3701 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3702 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3703 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3704 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3705 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3706 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3707 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3708 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3709 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3710 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3711 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3712 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3713 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3714 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3715 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3716 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3717 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3718 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3719 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3720 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3721 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3722 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3723 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3724 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3725 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3726 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3727 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3728 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3729 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3730 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3731 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3732 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3733 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3734 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3735 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3736 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3737 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3738 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3739 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3740 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3741 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3742 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3743 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3744 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3745 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3746 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3747 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3748 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3749 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3750 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3751 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3752 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3753 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3754 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3755 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3756 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3757 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3758 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3759 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3760 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3761 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3762 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3763 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3764 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3765 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3766 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3767 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3768 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3769 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3770 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3771 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3772 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3773 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3774 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3775 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3776 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3777 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3778 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3779 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3780 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3781 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3782 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3783 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3784 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3785 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3786 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3787 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3788 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3789 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3790 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3791 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3792 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3793 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3794 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3795 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3796 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3797 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3798 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3799 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3800 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3801 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3802 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3803 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3804 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3805 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3806 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3807 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3808 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3809 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3810 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3811 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3812 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3813 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3814 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3815 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3816 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3817 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3818 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3819 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3820 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3821 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3822 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3823 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3824 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3825 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3826 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3827 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3828 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3829 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3830 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3831 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3832 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3833 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3834 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3835 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3836 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3837 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3838 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3839 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3840 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3841 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3842 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3843 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3844 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3845 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3846 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3847 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3848 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3849 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3850 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3851 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3852 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3853 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3854 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3855 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3856 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3857 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3858 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3859 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3860 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3861 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3862 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3863 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3864 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3865 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3866 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3867 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3868 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3869 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3870 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3871 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3872 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3873 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3874 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3875 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3876 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3877 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3878 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3879 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3880 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3881 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3882 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3883 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3884 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3885 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3886 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3887 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3888 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3889 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3890 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3891 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3892 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3893 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3894 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3895 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3896 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3897 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3898 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3899 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3900 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3901 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3902 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3903 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3904 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3905 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3906 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3907 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3908 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3909 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3910 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3911 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3912 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3913 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3914 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3915 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3916 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3917 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3918 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3919 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3920 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3921 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3922 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3923 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3924 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3925 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3926 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3927 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3928 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3929 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3930 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3931 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3932 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3933 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3934 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3935 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3936 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3937 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3938 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3939 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3940 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3941 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3942 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3943 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3944 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3945 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3946 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3947 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3948 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3949 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3950 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3951 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3952 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3953 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3954 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3955 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3956 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3957 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3958 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3959 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3960 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3961 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3962 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3963 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3964 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3965 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3966 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3967 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3968 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3969 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3970 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3971 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3972 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3973 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3974 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3975 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3976 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3977 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3978 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3979 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3980 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3981 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3982 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3983 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3984 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3985 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3986 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3987 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3988 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3989 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3990 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3991 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3992 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3993 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3994 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3995 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3996 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3997 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3998 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3999 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4000 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4001 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4002 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4003 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4004 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4005 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4006 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4007 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4008 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4009 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4010 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4011 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4012 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4013 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4014 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4015 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4016 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4017 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4018 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4019 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4020 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4021 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4022 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4023 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4024 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4025 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4026 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4027 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4028 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4029 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4030 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4031 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4032 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4033 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4034 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4035 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4036 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4037 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4038 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4039 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4040 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4041 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4042 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4043 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4044 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4045 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4046 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4047 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4048 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4049 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4050 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4051 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4052 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4053 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4054 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4055 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4056 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4057 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4058 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4059 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4060 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4061 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4062 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4063 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4064 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4065 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4066 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4067 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4068 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4069 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4070 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4071 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4072 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4073 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4074 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4075 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4076 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4077 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4078 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4079 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4080 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4081 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4082 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4083 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4084 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4085 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4086 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4087 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4088 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4089 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4090 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4091 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4092 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4093 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4094 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4095 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4096 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4097 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4098 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4099 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4100 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4101 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4102 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4103 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4104 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4105 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4106 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4107 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4108 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4109 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4110 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4111 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4112 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4113 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4114 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4115 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4116 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4117 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4118 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4119 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4120 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4121 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4122 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4123 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4124 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4125 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4126 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4127 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4128 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4129 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4130 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4131 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4132 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4133 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4134 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4135 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4136 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4137 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4138 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4139 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4140 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4141 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4142 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4143 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4144 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4145 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4146 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4147 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4148 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4149 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4150 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4151 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4152 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4153 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4154 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4155 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4156 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4157 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4158 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4159 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4160 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4161 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4162 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4163 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4164 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4165 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4166 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4167 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4168 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4169 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4170 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4171 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4172 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4173 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4174 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4175 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4176 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4177 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4178 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4179 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4180 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4181 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4182 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4183 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4184 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4185 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4186 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4187 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4188 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4189 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4190 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4191 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4192 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4193 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4194 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4195 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4196 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4197 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4198 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4199 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4200 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4201 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4202 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4203 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4204 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4205 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4206 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4207 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4208 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4209 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4210 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4211 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4212 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4213 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4214 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4215 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4216 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4217 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4218 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4219 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4220 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4221 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4222 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4223 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4224 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4225 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4226 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4227 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4228 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4229 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4230 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4231 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4232 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4233 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4234 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4235 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4236 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4237 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4238 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4239 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4240 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4241 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4242 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4243 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4244 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4245 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4246 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4247 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4248 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4249 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4250 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4251 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4252 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4253 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4254 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4255 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4256 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4257 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4258 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4259 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4260 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4261 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4262 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4263 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4264 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4265 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4266 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4267 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4268 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4269 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4270 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4271 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4272 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4273 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4274 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4275 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4276 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4277 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4278 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4279 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4280 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4281 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4282 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4283 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4284 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4285 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4286 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4287 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4288 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4289 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4290 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4291 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4292 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4293 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4294 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4295 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4296 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4297 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4298 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4299 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4300 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4301 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4302 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4303 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4304 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4305 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4306 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4307 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4308 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4309 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4310 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4311 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4312 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4313 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4314 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4315 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4316 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4317 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4318 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4319 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4320 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4321 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4322 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4323 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4324 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4325 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4326 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4327 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4328 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4329 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4330 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4331 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4332 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4333 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4334 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4335 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4336 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4337 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4338 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4339 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4340 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4341 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4342 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4343 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4344 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4345 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4346 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4347 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4348 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4349 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4350 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4351 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4352 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4353 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4354 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4355 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4356 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4357 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4358 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4359 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4360 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4361 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4362 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4363 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4364 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4365 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4366 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4367 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4368 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4369 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4370 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4371 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4372 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4373 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4374 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4375 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4376 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4377 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4378 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4379 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4380 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4381 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4382 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4383 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4384 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4385 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4386 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4387 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4388 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4389 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4390 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4391 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4392 outd_stage2_3/cmirror_out m2_40400_10380# m4_40470_12880# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4393 m4_40470_12880# m2_40400_10380# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4394 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4395 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4396 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4397 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4398 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4399 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4400 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4401 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4402 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4403 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4404 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4405 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4406 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4407 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4408 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4409 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4410 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4411 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4412 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4413 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4414 outd_stage2_3/cmirror_out m2_40400_9110# m4_40470_12200# outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4415 m4_40470_12200# m2_40400_9110# outd_stage2_3/cmirror_out outd_stage2_3/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4416 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4417 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4418 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4419 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4420 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4421 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4422 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4423 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4424 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4425 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4426 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4427 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4428 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4429 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4430 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4431 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4432 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4433 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4434 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4435 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4436 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4437 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4438 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4439 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4440 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4441 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4442 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4443 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4444 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4445 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4446 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4447 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4448 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4449 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4450 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4451 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4452 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4453 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4454 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4455 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4456 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4457 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4458 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4459 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4460 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4461 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4462 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4463 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4464 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4465 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4466 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4467 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4468 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4469 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4470 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4471 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4472 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4473 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4474 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4475 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4476 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4477 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4478 outd_stage2_3/cmirror_out outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4479 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# outd_stage2_3/cmirror_out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4480 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4481 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4482 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4483 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4484 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4485 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4486 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4487 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4488 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4489 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4490 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4491 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4492 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4493 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4494 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4495 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4496 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4497 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4498 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4499 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4500 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4501 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4502 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4503 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4504 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4505 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4506 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4507 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4508 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4509 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4510 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4511 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4512 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4513 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4514 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4515 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4516 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4517 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4518 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4519 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4520 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4521 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4522 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4523 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4524 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4525 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4526 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4527 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4528 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4529 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4530 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4531 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4532 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4533 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4534 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4535 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4536 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4537 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4538 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4539 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4540 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4541 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4542 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4543 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4544 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4545 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4546 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4547 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4548 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4549 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4550 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4551 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4552 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4553 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4554 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4555 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4556 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4557 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4558 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4559 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4560 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4561 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4562 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4563 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4564 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4565 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4566 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4567 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4568 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4569 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4570 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4571 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4572 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4573 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4574 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4575 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4576 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4577 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4578 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4579 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4580 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4581 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4582 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4583 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4584 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4585 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4586 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4587 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4588 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4589 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4590 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4591 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4592 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4593 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4594 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4595 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4596 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4597 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4598 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4599 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4600 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4601 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4602 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4603 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4604 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4605 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4606 VSUBS outd_stage2_3/outd_cmirror_64t_4/m1_0_80# m2_41490_8160# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4607 m2_41490_8160# outd_stage2_3/outd_cmirror_64t_4/m1_0_80# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
