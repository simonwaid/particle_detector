magic
tech sky130A
magscale 1 2
timestamp 1645781187
<< error_p >>
rect -715 581 -657 587
rect -519 581 -461 587
rect -323 581 -265 587
rect -127 581 -69 587
rect 69 581 127 587
rect 265 581 323 587
rect 461 581 519 587
rect 657 581 715 587
rect -715 547 -703 581
rect -519 547 -507 581
rect -323 547 -311 581
rect -127 547 -115 581
rect 69 547 81 581
rect 265 547 277 581
rect 461 547 473 581
rect 657 547 669 581
rect -715 541 -657 547
rect -519 541 -461 547
rect -323 541 -265 547
rect -127 541 -69 547
rect 69 541 127 547
rect 265 541 323 547
rect 461 541 519 547
rect 657 541 715 547
rect -617 71 -559 77
rect -421 71 -363 77
rect -225 71 -167 77
rect -29 71 29 77
rect 167 71 225 77
rect 363 71 421 77
rect 559 71 617 77
rect -617 37 -605 71
rect -421 37 -409 71
rect -225 37 -213 71
rect -29 37 -17 71
rect 167 37 179 71
rect 363 37 375 71
rect 559 37 571 71
rect -617 31 -559 37
rect -421 31 -363 37
rect -225 31 -167 37
rect -29 31 29 37
rect 167 31 225 37
rect 363 31 421 37
rect 559 31 617 37
rect -617 -37 -559 -31
rect -421 -37 -363 -31
rect -225 -37 -167 -31
rect -29 -37 29 -31
rect 167 -37 225 -31
rect 363 -37 421 -31
rect 559 -37 617 -31
rect -617 -71 -605 -37
rect -421 -71 -409 -37
rect -225 -71 -213 -37
rect -29 -71 -17 -37
rect 167 -71 179 -37
rect 363 -71 375 -37
rect 559 -71 571 -37
rect -617 -77 -559 -71
rect -421 -77 -363 -71
rect -225 -77 -167 -71
rect -29 -77 29 -71
rect 167 -77 225 -71
rect 363 -77 421 -71
rect 559 -77 617 -71
rect -715 -547 -657 -541
rect -519 -547 -461 -541
rect -323 -547 -265 -541
rect -127 -547 -69 -541
rect 69 -547 127 -541
rect 265 -547 323 -541
rect 461 -547 519 -541
rect 657 -547 715 -541
rect -715 -581 -703 -547
rect -519 -581 -507 -547
rect -323 -581 -311 -547
rect -127 -581 -115 -547
rect 69 -581 81 -547
rect 265 -581 277 -547
rect 461 -581 473 -547
rect 657 -581 669 -547
rect -715 -587 -657 -581
rect -519 -587 -461 -581
rect -323 -587 -265 -581
rect -127 -587 -69 -581
rect 69 -587 127 -581
rect 265 -587 323 -581
rect 461 -587 519 -581
rect 657 -587 715 -581
<< pwell >>
rect -902 -719 902 719
<< nmos >>
rect -706 109 -666 509
rect -608 109 -568 509
rect -510 109 -470 509
rect -412 109 -372 509
rect -314 109 -274 509
rect -216 109 -176 509
rect -118 109 -78 509
rect -20 109 20 509
rect 78 109 118 509
rect 176 109 216 509
rect 274 109 314 509
rect 372 109 412 509
rect 470 109 510 509
rect 568 109 608 509
rect 666 109 706 509
rect -706 -509 -666 -109
rect -608 -509 -568 -109
rect -510 -509 -470 -109
rect -412 -509 -372 -109
rect -314 -509 -274 -109
rect -216 -509 -176 -109
rect -118 -509 -78 -109
rect -20 -509 20 -109
rect 78 -509 118 -109
rect 176 -509 216 -109
rect 274 -509 314 -109
rect 372 -509 412 -109
rect 470 -509 510 -109
rect 568 -509 608 -109
rect 666 -509 706 -109
<< ndiff >>
rect -764 497 -706 509
rect -764 121 -752 497
rect -718 121 -706 497
rect -764 109 -706 121
rect -666 497 -608 509
rect -666 121 -654 497
rect -620 121 -608 497
rect -666 109 -608 121
rect -568 497 -510 509
rect -568 121 -556 497
rect -522 121 -510 497
rect -568 109 -510 121
rect -470 497 -412 509
rect -470 121 -458 497
rect -424 121 -412 497
rect -470 109 -412 121
rect -372 497 -314 509
rect -372 121 -360 497
rect -326 121 -314 497
rect -372 109 -314 121
rect -274 497 -216 509
rect -274 121 -262 497
rect -228 121 -216 497
rect -274 109 -216 121
rect -176 497 -118 509
rect -176 121 -164 497
rect -130 121 -118 497
rect -176 109 -118 121
rect -78 497 -20 509
rect -78 121 -66 497
rect -32 121 -20 497
rect -78 109 -20 121
rect 20 497 78 509
rect 20 121 32 497
rect 66 121 78 497
rect 20 109 78 121
rect 118 497 176 509
rect 118 121 130 497
rect 164 121 176 497
rect 118 109 176 121
rect 216 497 274 509
rect 216 121 228 497
rect 262 121 274 497
rect 216 109 274 121
rect 314 497 372 509
rect 314 121 326 497
rect 360 121 372 497
rect 314 109 372 121
rect 412 497 470 509
rect 412 121 424 497
rect 458 121 470 497
rect 412 109 470 121
rect 510 497 568 509
rect 510 121 522 497
rect 556 121 568 497
rect 510 109 568 121
rect 608 497 666 509
rect 608 121 620 497
rect 654 121 666 497
rect 608 109 666 121
rect 706 497 764 509
rect 706 121 718 497
rect 752 121 764 497
rect 706 109 764 121
rect -764 -121 -706 -109
rect -764 -497 -752 -121
rect -718 -497 -706 -121
rect -764 -509 -706 -497
rect -666 -121 -608 -109
rect -666 -497 -654 -121
rect -620 -497 -608 -121
rect -666 -509 -608 -497
rect -568 -121 -510 -109
rect -568 -497 -556 -121
rect -522 -497 -510 -121
rect -568 -509 -510 -497
rect -470 -121 -412 -109
rect -470 -497 -458 -121
rect -424 -497 -412 -121
rect -470 -509 -412 -497
rect -372 -121 -314 -109
rect -372 -497 -360 -121
rect -326 -497 -314 -121
rect -372 -509 -314 -497
rect -274 -121 -216 -109
rect -274 -497 -262 -121
rect -228 -497 -216 -121
rect -274 -509 -216 -497
rect -176 -121 -118 -109
rect -176 -497 -164 -121
rect -130 -497 -118 -121
rect -176 -509 -118 -497
rect -78 -121 -20 -109
rect -78 -497 -66 -121
rect -32 -497 -20 -121
rect -78 -509 -20 -497
rect 20 -121 78 -109
rect 20 -497 32 -121
rect 66 -497 78 -121
rect 20 -509 78 -497
rect 118 -121 176 -109
rect 118 -497 130 -121
rect 164 -497 176 -121
rect 118 -509 176 -497
rect 216 -121 274 -109
rect 216 -497 228 -121
rect 262 -497 274 -121
rect 216 -509 274 -497
rect 314 -121 372 -109
rect 314 -497 326 -121
rect 360 -497 372 -121
rect 314 -509 372 -497
rect 412 -121 470 -109
rect 412 -497 424 -121
rect 458 -497 470 -121
rect 412 -509 470 -497
rect 510 -121 568 -109
rect 510 -497 522 -121
rect 556 -497 568 -121
rect 510 -509 568 -497
rect 608 -121 666 -109
rect 608 -497 620 -121
rect 654 -497 666 -121
rect 608 -509 666 -497
rect 706 -121 764 -109
rect 706 -497 718 -121
rect 752 -497 764 -121
rect 706 -509 764 -497
<< ndiffc >>
rect -752 121 -718 497
rect -654 121 -620 497
rect -556 121 -522 497
rect -458 121 -424 497
rect -360 121 -326 497
rect -262 121 -228 497
rect -164 121 -130 497
rect -66 121 -32 497
rect 32 121 66 497
rect 130 121 164 497
rect 228 121 262 497
rect 326 121 360 497
rect 424 121 458 497
rect 522 121 556 497
rect 620 121 654 497
rect 718 121 752 497
rect -752 -497 -718 -121
rect -654 -497 -620 -121
rect -556 -497 -522 -121
rect -458 -497 -424 -121
rect -360 -497 -326 -121
rect -262 -497 -228 -121
rect -164 -497 -130 -121
rect -66 -497 -32 -121
rect 32 -497 66 -121
rect 130 -497 164 -121
rect 228 -497 262 -121
rect 326 -497 360 -121
rect 424 -497 458 -121
rect 522 -497 556 -121
rect 620 -497 654 -121
rect 718 -497 752 -121
<< psubdiff >>
rect -866 649 -770 683
rect 770 649 866 683
rect -866 587 -832 649
rect 832 587 866 649
rect -866 -649 -832 -587
rect 832 -649 866 -587
rect -866 -683 -770 -649
rect 770 -683 866 -649
<< psubdiffcont >>
rect -770 649 770 683
rect -866 -587 -832 587
rect 832 -587 866 587
rect -770 -683 770 -649
<< poly >>
rect -719 581 -653 597
rect -719 547 -703 581
rect -669 547 -653 581
rect -719 531 -653 547
rect -523 581 -457 597
rect -523 547 -507 581
rect -473 547 -457 581
rect -706 509 -666 531
rect -608 509 -568 535
rect -523 531 -457 547
rect -327 581 -261 597
rect -327 547 -311 581
rect -277 547 -261 581
rect -510 509 -470 531
rect -412 509 -372 535
rect -327 531 -261 547
rect -131 581 -65 597
rect -131 547 -115 581
rect -81 547 -65 581
rect -314 509 -274 531
rect -216 509 -176 535
rect -131 531 -65 547
rect 65 581 131 597
rect 65 547 81 581
rect 115 547 131 581
rect -118 509 -78 531
rect -20 509 20 535
rect 65 531 131 547
rect 261 581 327 597
rect 261 547 277 581
rect 311 547 327 581
rect 78 509 118 531
rect 176 509 216 535
rect 261 531 327 547
rect 457 581 523 597
rect 457 547 473 581
rect 507 547 523 581
rect 274 509 314 531
rect 372 509 412 535
rect 457 531 523 547
rect 653 581 719 597
rect 653 547 669 581
rect 703 547 719 581
rect 470 509 510 531
rect 568 509 608 535
rect 653 531 719 547
rect 666 509 706 531
rect -706 83 -666 109
rect -608 87 -568 109
rect -621 71 -555 87
rect -510 83 -470 109
rect -412 87 -372 109
rect -621 37 -605 71
rect -571 37 -555 71
rect -621 21 -555 37
rect -425 71 -359 87
rect -314 83 -274 109
rect -216 87 -176 109
rect -425 37 -409 71
rect -375 37 -359 71
rect -425 21 -359 37
rect -229 71 -163 87
rect -118 83 -78 109
rect -20 87 20 109
rect -229 37 -213 71
rect -179 37 -163 71
rect -229 21 -163 37
rect -33 71 33 87
rect 78 83 118 109
rect 176 87 216 109
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 163 71 229 87
rect 274 83 314 109
rect 372 87 412 109
rect 163 37 179 71
rect 213 37 229 71
rect 163 21 229 37
rect 359 71 425 87
rect 470 83 510 109
rect 568 87 608 109
rect 359 37 375 71
rect 409 37 425 71
rect 359 21 425 37
rect 555 71 621 87
rect 666 83 706 109
rect 555 37 571 71
rect 605 37 621 71
rect 555 21 621 37
rect -621 -37 -555 -21
rect -621 -71 -605 -37
rect -571 -71 -555 -37
rect -706 -109 -666 -83
rect -621 -87 -555 -71
rect -425 -37 -359 -21
rect -425 -71 -409 -37
rect -375 -71 -359 -37
rect -608 -109 -568 -87
rect -510 -109 -470 -83
rect -425 -87 -359 -71
rect -229 -37 -163 -21
rect -229 -71 -213 -37
rect -179 -71 -163 -37
rect -412 -109 -372 -87
rect -314 -109 -274 -83
rect -229 -87 -163 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -216 -109 -176 -87
rect -118 -109 -78 -83
rect -33 -87 33 -71
rect 163 -37 229 -21
rect 163 -71 179 -37
rect 213 -71 229 -37
rect -20 -109 20 -87
rect 78 -109 118 -83
rect 163 -87 229 -71
rect 359 -37 425 -21
rect 359 -71 375 -37
rect 409 -71 425 -37
rect 176 -109 216 -87
rect 274 -109 314 -83
rect 359 -87 425 -71
rect 555 -37 621 -21
rect 555 -71 571 -37
rect 605 -71 621 -37
rect 372 -109 412 -87
rect 470 -109 510 -83
rect 555 -87 621 -71
rect 568 -109 608 -87
rect 666 -109 706 -83
rect -706 -531 -666 -509
rect -719 -547 -653 -531
rect -608 -535 -568 -509
rect -510 -531 -470 -509
rect -719 -581 -703 -547
rect -669 -581 -653 -547
rect -719 -597 -653 -581
rect -523 -547 -457 -531
rect -412 -535 -372 -509
rect -314 -531 -274 -509
rect -523 -581 -507 -547
rect -473 -581 -457 -547
rect -523 -597 -457 -581
rect -327 -547 -261 -531
rect -216 -535 -176 -509
rect -118 -531 -78 -509
rect -327 -581 -311 -547
rect -277 -581 -261 -547
rect -327 -597 -261 -581
rect -131 -547 -65 -531
rect -20 -535 20 -509
rect 78 -531 118 -509
rect -131 -581 -115 -547
rect -81 -581 -65 -547
rect -131 -597 -65 -581
rect 65 -547 131 -531
rect 176 -535 216 -509
rect 274 -531 314 -509
rect 65 -581 81 -547
rect 115 -581 131 -547
rect 65 -597 131 -581
rect 261 -547 327 -531
rect 372 -535 412 -509
rect 470 -531 510 -509
rect 261 -581 277 -547
rect 311 -581 327 -547
rect 261 -597 327 -581
rect 457 -547 523 -531
rect 568 -535 608 -509
rect 666 -531 706 -509
rect 457 -581 473 -547
rect 507 -581 523 -547
rect 457 -597 523 -581
rect 653 -547 719 -531
rect 653 -581 669 -547
rect 703 -581 719 -547
rect 653 -597 719 -581
<< polycont >>
rect -703 547 -669 581
rect -507 547 -473 581
rect -311 547 -277 581
rect -115 547 -81 581
rect 81 547 115 581
rect 277 547 311 581
rect 473 547 507 581
rect 669 547 703 581
rect -605 37 -571 71
rect -409 37 -375 71
rect -213 37 -179 71
rect -17 37 17 71
rect 179 37 213 71
rect 375 37 409 71
rect 571 37 605 71
rect -605 -71 -571 -37
rect -409 -71 -375 -37
rect -213 -71 -179 -37
rect -17 -71 17 -37
rect 179 -71 213 -37
rect 375 -71 409 -37
rect 571 -71 605 -37
rect -703 -581 -669 -547
rect -507 -581 -473 -547
rect -311 -581 -277 -547
rect -115 -581 -81 -547
rect 81 -581 115 -547
rect 277 -581 311 -547
rect 473 -581 507 -547
rect 669 -581 703 -547
<< locali >>
rect -866 649 -770 683
rect 770 649 866 683
rect -866 587 -832 649
rect 832 587 866 649
rect -719 547 -703 581
rect -669 547 -653 581
rect -523 547 -507 581
rect -473 547 -457 581
rect -327 547 -311 581
rect -277 547 -261 581
rect -131 547 -115 581
rect -81 547 -65 581
rect 65 547 81 581
rect 115 547 131 581
rect 261 547 277 581
rect 311 547 327 581
rect 457 547 473 581
rect 507 547 523 581
rect 653 547 669 581
rect 703 547 719 581
rect -752 497 -718 513
rect -752 105 -718 121
rect -654 497 -620 513
rect -654 105 -620 121
rect -556 497 -522 513
rect -556 105 -522 121
rect -458 497 -424 513
rect -458 105 -424 121
rect -360 497 -326 513
rect -360 105 -326 121
rect -262 497 -228 513
rect -262 105 -228 121
rect -164 497 -130 513
rect -164 105 -130 121
rect -66 497 -32 513
rect -66 105 -32 121
rect 32 497 66 513
rect 32 105 66 121
rect 130 497 164 513
rect 130 105 164 121
rect 228 497 262 513
rect 228 105 262 121
rect 326 497 360 513
rect 326 105 360 121
rect 424 497 458 513
rect 424 105 458 121
rect 522 497 556 513
rect 522 105 556 121
rect 620 497 654 513
rect 620 105 654 121
rect 718 497 752 513
rect 718 105 752 121
rect -621 37 -605 71
rect -571 37 -555 71
rect -425 37 -409 71
rect -375 37 -359 71
rect -229 37 -213 71
rect -179 37 -163 71
rect -33 37 -17 71
rect 17 37 33 71
rect 163 37 179 71
rect 213 37 229 71
rect 359 37 375 71
rect 409 37 425 71
rect 555 37 571 71
rect 605 37 621 71
rect -621 -71 -605 -37
rect -571 -71 -555 -37
rect -425 -71 -409 -37
rect -375 -71 -359 -37
rect -229 -71 -213 -37
rect -179 -71 -163 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 163 -71 179 -37
rect 213 -71 229 -37
rect 359 -71 375 -37
rect 409 -71 425 -37
rect 555 -71 571 -37
rect 605 -71 621 -37
rect -752 -121 -718 -105
rect -752 -513 -718 -497
rect -654 -121 -620 -105
rect -654 -513 -620 -497
rect -556 -121 -522 -105
rect -556 -513 -522 -497
rect -458 -121 -424 -105
rect -458 -513 -424 -497
rect -360 -121 -326 -105
rect -360 -513 -326 -497
rect -262 -121 -228 -105
rect -262 -513 -228 -497
rect -164 -121 -130 -105
rect -164 -513 -130 -497
rect -66 -121 -32 -105
rect -66 -513 -32 -497
rect 32 -121 66 -105
rect 32 -513 66 -497
rect 130 -121 164 -105
rect 130 -513 164 -497
rect 228 -121 262 -105
rect 228 -513 262 -497
rect 326 -121 360 -105
rect 326 -513 360 -497
rect 424 -121 458 -105
rect 424 -513 458 -497
rect 522 -121 556 -105
rect 522 -513 556 -497
rect 620 -121 654 -105
rect 620 -513 654 -497
rect 718 -121 752 -105
rect 718 -513 752 -497
rect -719 -581 -703 -547
rect -669 -581 -653 -547
rect -523 -581 -507 -547
rect -473 -581 -457 -547
rect -327 -581 -311 -547
rect -277 -581 -261 -547
rect -131 -581 -115 -547
rect -81 -581 -65 -547
rect 65 -581 81 -547
rect 115 -581 131 -547
rect 261 -581 277 -547
rect 311 -581 327 -547
rect 457 -581 473 -547
rect 507 -581 523 -547
rect 653 -581 669 -547
rect 703 -581 719 -547
rect -866 -649 -832 -587
rect 832 -649 866 -587
rect -866 -683 -770 -649
rect 770 -683 866 -649
<< viali >>
rect -703 547 -669 581
rect -507 547 -473 581
rect -311 547 -277 581
rect -115 547 -81 581
rect 81 547 115 581
rect 277 547 311 581
rect 473 547 507 581
rect 669 547 703 581
rect -752 121 -718 497
rect -654 121 -620 497
rect -556 121 -522 497
rect -458 121 -424 497
rect -360 121 -326 497
rect -262 121 -228 497
rect -164 121 -130 497
rect -66 121 -32 497
rect 32 121 66 497
rect 130 121 164 497
rect 228 121 262 497
rect 326 121 360 497
rect 424 121 458 497
rect 522 121 556 497
rect 620 121 654 497
rect 718 121 752 497
rect -605 37 -571 71
rect -409 37 -375 71
rect -213 37 -179 71
rect -17 37 17 71
rect 179 37 213 71
rect 375 37 409 71
rect 571 37 605 71
rect -605 -71 -571 -37
rect -409 -71 -375 -37
rect -213 -71 -179 -37
rect -17 -71 17 -37
rect 179 -71 213 -37
rect 375 -71 409 -37
rect 571 -71 605 -37
rect -752 -497 -718 -121
rect -654 -497 -620 -121
rect -556 -497 -522 -121
rect -458 -497 -424 -121
rect -360 -497 -326 -121
rect -262 -497 -228 -121
rect -164 -497 -130 -121
rect -66 -497 -32 -121
rect 32 -497 66 -121
rect 130 -497 164 -121
rect 228 -497 262 -121
rect 326 -497 360 -121
rect 424 -497 458 -121
rect 522 -497 556 -121
rect 620 -497 654 -121
rect 718 -497 752 -121
rect -703 -581 -669 -547
rect -507 -581 -473 -547
rect -311 -581 -277 -547
rect -115 -581 -81 -547
rect 81 -581 115 -547
rect 277 -581 311 -547
rect 473 -581 507 -547
rect 669 -581 703 -547
<< metal1 >>
rect -715 581 -657 587
rect -715 547 -703 581
rect -669 547 -657 581
rect -715 541 -657 547
rect -519 581 -461 587
rect -519 547 -507 581
rect -473 547 -461 581
rect -519 541 -461 547
rect -323 581 -265 587
rect -323 547 -311 581
rect -277 547 -265 581
rect -323 541 -265 547
rect -127 581 -69 587
rect -127 547 -115 581
rect -81 547 -69 581
rect -127 541 -69 547
rect 69 581 127 587
rect 69 547 81 581
rect 115 547 127 581
rect 69 541 127 547
rect 265 581 323 587
rect 265 547 277 581
rect 311 547 323 581
rect 265 541 323 547
rect 461 581 519 587
rect 461 547 473 581
rect 507 547 519 581
rect 461 541 519 547
rect 657 581 715 587
rect 657 547 669 581
rect 703 547 715 581
rect 657 541 715 547
rect -758 497 -712 509
rect -758 121 -752 497
rect -718 121 -712 497
rect -758 109 -712 121
rect -660 497 -614 509
rect -660 121 -654 497
rect -620 121 -614 497
rect -660 109 -614 121
rect -562 497 -516 509
rect -562 121 -556 497
rect -522 121 -516 497
rect -562 109 -516 121
rect -464 497 -418 509
rect -464 121 -458 497
rect -424 121 -418 497
rect -464 109 -418 121
rect -366 497 -320 509
rect -366 121 -360 497
rect -326 121 -320 497
rect -366 109 -320 121
rect -268 497 -222 509
rect -268 121 -262 497
rect -228 121 -222 497
rect -268 109 -222 121
rect -170 497 -124 509
rect -170 121 -164 497
rect -130 121 -124 497
rect -170 109 -124 121
rect -72 497 -26 509
rect -72 121 -66 497
rect -32 121 -26 497
rect -72 109 -26 121
rect 26 497 72 509
rect 26 121 32 497
rect 66 121 72 497
rect 26 109 72 121
rect 124 497 170 509
rect 124 121 130 497
rect 164 121 170 497
rect 124 109 170 121
rect 222 497 268 509
rect 222 121 228 497
rect 262 121 268 497
rect 222 109 268 121
rect 320 497 366 509
rect 320 121 326 497
rect 360 121 366 497
rect 320 109 366 121
rect 418 497 464 509
rect 418 121 424 497
rect 458 121 464 497
rect 418 109 464 121
rect 516 497 562 509
rect 516 121 522 497
rect 556 121 562 497
rect 516 109 562 121
rect 614 497 660 509
rect 614 121 620 497
rect 654 121 660 497
rect 614 109 660 121
rect 712 497 758 509
rect 712 121 718 497
rect 752 121 758 497
rect 712 109 758 121
rect -617 71 -559 77
rect -617 37 -605 71
rect -571 37 -559 71
rect -617 31 -559 37
rect -421 71 -363 77
rect -421 37 -409 71
rect -375 37 -363 71
rect -421 31 -363 37
rect -225 71 -167 77
rect -225 37 -213 71
rect -179 37 -167 71
rect -225 31 -167 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 167 71 225 77
rect 167 37 179 71
rect 213 37 225 71
rect 167 31 225 37
rect 363 71 421 77
rect 363 37 375 71
rect 409 37 421 71
rect 363 31 421 37
rect 559 71 617 77
rect 559 37 571 71
rect 605 37 617 71
rect 559 31 617 37
rect -617 -37 -559 -31
rect -617 -71 -605 -37
rect -571 -71 -559 -37
rect -617 -77 -559 -71
rect -421 -37 -363 -31
rect -421 -71 -409 -37
rect -375 -71 -363 -37
rect -421 -77 -363 -71
rect -225 -37 -167 -31
rect -225 -71 -213 -37
rect -179 -71 -167 -37
rect -225 -77 -167 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 167 -37 225 -31
rect 167 -71 179 -37
rect 213 -71 225 -37
rect 167 -77 225 -71
rect 363 -37 421 -31
rect 363 -71 375 -37
rect 409 -71 421 -37
rect 363 -77 421 -71
rect 559 -37 617 -31
rect 559 -71 571 -37
rect 605 -71 617 -37
rect 559 -77 617 -71
rect -758 -121 -712 -109
rect -758 -497 -752 -121
rect -718 -497 -712 -121
rect -758 -509 -712 -497
rect -660 -121 -614 -109
rect -660 -497 -654 -121
rect -620 -497 -614 -121
rect -660 -509 -614 -497
rect -562 -121 -516 -109
rect -562 -497 -556 -121
rect -522 -497 -516 -121
rect -562 -509 -516 -497
rect -464 -121 -418 -109
rect -464 -497 -458 -121
rect -424 -497 -418 -121
rect -464 -509 -418 -497
rect -366 -121 -320 -109
rect -366 -497 -360 -121
rect -326 -497 -320 -121
rect -366 -509 -320 -497
rect -268 -121 -222 -109
rect -268 -497 -262 -121
rect -228 -497 -222 -121
rect -268 -509 -222 -497
rect -170 -121 -124 -109
rect -170 -497 -164 -121
rect -130 -497 -124 -121
rect -170 -509 -124 -497
rect -72 -121 -26 -109
rect -72 -497 -66 -121
rect -32 -497 -26 -121
rect -72 -509 -26 -497
rect 26 -121 72 -109
rect 26 -497 32 -121
rect 66 -497 72 -121
rect 26 -509 72 -497
rect 124 -121 170 -109
rect 124 -497 130 -121
rect 164 -497 170 -121
rect 124 -509 170 -497
rect 222 -121 268 -109
rect 222 -497 228 -121
rect 262 -497 268 -121
rect 222 -509 268 -497
rect 320 -121 366 -109
rect 320 -497 326 -121
rect 360 -497 366 -121
rect 320 -509 366 -497
rect 418 -121 464 -109
rect 418 -497 424 -121
rect 458 -497 464 -121
rect 418 -509 464 -497
rect 516 -121 562 -109
rect 516 -497 522 -121
rect 556 -497 562 -121
rect 516 -509 562 -497
rect 614 -121 660 -109
rect 614 -497 620 -121
rect 654 -497 660 -121
rect 614 -509 660 -497
rect 712 -121 758 -109
rect 712 -497 718 -121
rect 752 -497 758 -121
rect 712 -509 758 -497
rect -715 -547 -657 -541
rect -715 -581 -703 -547
rect -669 -581 -657 -547
rect -715 -587 -657 -581
rect -519 -547 -461 -541
rect -519 -581 -507 -547
rect -473 -581 -461 -547
rect -519 -587 -461 -581
rect -323 -547 -265 -541
rect -323 -581 -311 -547
rect -277 -581 -265 -547
rect -323 -587 -265 -581
rect -127 -547 -69 -541
rect -127 -581 -115 -547
rect -81 -581 -69 -547
rect -127 -587 -69 -581
rect 69 -547 127 -541
rect 69 -581 81 -547
rect 115 -581 127 -547
rect 69 -587 127 -581
rect 265 -547 323 -541
rect 265 -581 277 -547
rect 311 -581 323 -547
rect 265 -587 323 -581
rect 461 -547 519 -541
rect 461 -581 473 -547
rect 507 -581 519 -547
rect 461 -587 519 -581
rect 657 -547 715 -541
rect 657 -581 669 -547
rect 703 -581 715 -547
rect 657 -587 715 -581
<< properties >>
string FIXED_BBOX -849 -666 849 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.2 m 2 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
