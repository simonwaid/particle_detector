magic
tech sky130A
magscale 1 2
timestamp 1646400034
<< nwell >>
rect -1883 -319 1883 319
<< pmos >>
rect -1687 -100 -887 100
rect -829 -100 -29 100
rect 29 -100 829 100
rect 887 -100 1687 100
<< pdiff >>
rect -1745 88 -1687 100
rect -1745 -88 -1733 88
rect -1699 -88 -1687 88
rect -1745 -100 -1687 -88
rect -887 88 -829 100
rect -887 -88 -875 88
rect -841 -88 -829 88
rect -887 -100 -829 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 829 88 887 100
rect 829 -88 841 88
rect 875 -88 887 88
rect 829 -100 887 -88
rect 1687 88 1745 100
rect 1687 -88 1699 88
rect 1733 -88 1745 88
rect 1687 -100 1745 -88
<< pdiffc >>
rect -1733 -88 -1699 88
rect -875 -88 -841 88
rect -17 -88 17 88
rect 841 -88 875 88
rect 1699 -88 1733 88
<< nsubdiff >>
rect -1847 249 -1751 283
rect 1751 249 1847 283
rect -1847 187 -1813 249
rect 1813 187 1847 249
rect -1847 -249 -1813 -187
rect 1813 -249 1847 -187
rect -1847 -283 -1751 -249
rect 1751 -283 1847 -249
<< nsubdiffcont >>
rect -1751 249 1751 283
rect -1847 -187 -1813 187
rect 1813 -187 1847 187
rect -1751 -283 1751 -249
<< poly >>
rect -1687 181 -887 197
rect -1687 147 -1671 181
rect -903 147 -887 181
rect -1687 100 -887 147
rect -829 181 -29 197
rect -829 147 -813 181
rect -45 147 -29 181
rect -829 100 -29 147
rect 29 181 829 197
rect 29 147 45 181
rect 813 147 829 181
rect 29 100 829 147
rect 887 181 1687 197
rect 887 147 903 181
rect 1671 147 1687 181
rect 887 100 1687 147
rect -1687 -147 -887 -100
rect -1687 -181 -1671 -147
rect -903 -181 -887 -147
rect -1687 -197 -887 -181
rect -829 -147 -29 -100
rect -829 -181 -813 -147
rect -45 -181 -29 -147
rect -829 -197 -29 -181
rect 29 -147 829 -100
rect 29 -181 45 -147
rect 813 -181 829 -147
rect 29 -197 829 -181
rect 887 -147 1687 -100
rect 887 -181 903 -147
rect 1671 -181 1687 -147
rect 887 -197 1687 -181
<< polycont >>
rect -1671 147 -903 181
rect -813 147 -45 181
rect 45 147 813 181
rect 903 147 1671 181
rect -1671 -181 -903 -147
rect -813 -181 -45 -147
rect 45 -181 813 -147
rect 903 -181 1671 -147
<< locali >>
rect -1847 249 -1751 283
rect 1751 249 1847 283
rect -1847 187 -1813 249
rect 1813 187 1847 249
rect -1687 147 -1671 181
rect -903 147 -887 181
rect -829 147 -813 181
rect -45 147 -29 181
rect 29 147 45 181
rect 813 147 829 181
rect 887 147 903 181
rect 1671 147 1687 181
rect -1733 88 -1699 104
rect -1733 -104 -1699 -88
rect -875 88 -841 104
rect -875 -104 -841 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 841 88 875 104
rect 841 -104 875 -88
rect 1699 88 1733 104
rect 1699 -104 1733 -88
rect -1687 -181 -1671 -147
rect -903 -181 -887 -147
rect -829 -181 -813 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 813 -181 829 -147
rect 887 -181 903 -147
rect 1671 -181 1687 -147
rect -1847 -249 -1813 -187
rect 1813 -249 1847 -187
rect -1847 -283 -1751 -249
rect 1751 -283 1847 -249
<< viali >>
rect -1671 147 -903 181
rect -813 147 -45 181
rect 45 147 813 181
rect 903 147 1671 181
rect -1733 -88 -1699 88
rect -875 -88 -841 88
rect -17 -88 17 88
rect 841 -88 875 88
rect 1699 -88 1733 88
rect -1671 -181 -903 -147
rect -813 -181 -45 -147
rect 45 -181 813 -147
rect 903 -181 1671 -147
<< metal1 >>
rect -1683 181 -891 187
rect -1683 147 -1671 181
rect -903 147 -891 181
rect -1683 141 -891 147
rect -825 181 -33 187
rect -825 147 -813 181
rect -45 147 -33 181
rect -825 141 -33 147
rect 33 181 825 187
rect 33 147 45 181
rect 813 147 825 181
rect 33 141 825 147
rect 891 181 1683 187
rect 891 147 903 181
rect 1671 147 1683 181
rect 891 141 1683 147
rect -1739 88 -1693 100
rect -1739 -88 -1733 88
rect -1699 -88 -1693 88
rect -1739 -100 -1693 -88
rect -881 88 -835 100
rect -881 -88 -875 88
rect -841 -88 -835 88
rect -881 -100 -835 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 835 88 881 100
rect 835 -88 841 88
rect 875 -88 881 88
rect 835 -100 881 -88
rect 1693 88 1739 100
rect 1693 -88 1699 88
rect 1733 -88 1739 88
rect 1693 -100 1739 -88
rect -1683 -147 -891 -141
rect -1683 -181 -1671 -147
rect -903 -181 -891 -147
rect -1683 -187 -891 -181
rect -825 -147 -33 -141
rect -825 -181 -813 -147
rect -45 -181 -33 -147
rect -825 -187 -33 -181
rect 33 -147 825 -141
rect 33 -181 45 -147
rect 813 -181 825 -147
rect 33 -187 825 -181
rect 891 -147 1683 -141
rect 891 -181 903 -147
rect 1671 -181 1683 -147
rect 891 -187 1683 -181
<< properties >>
string FIXED_BBOX -1830 -266 1830 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 4 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
