** sch_path: /home/simon/code/caravel_tia/xschem/esd/esd_diodes.sch
**.subckt esd_diodes VP io VN
*.iopin VP
*.iopin io
*.iopin VN
D1 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D11 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D2 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D3 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D4 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D5 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D6 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D7 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D8 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D9 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D10 io VP sky130_fd_pr__diode_pd2nw_11v0 area=4e12
D12 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D13 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D14 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D15 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D16 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D17 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D18 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D19 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
D20 VN io sky130_fd_pr__diode_pw2nd_11v0 area=4e12
**.ends
.end
