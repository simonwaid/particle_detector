magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< error_p >>
rect -365 599 -307 605
rect -173 599 -115 605
rect 19 599 77 605
rect 211 599 269 605
rect -365 565 -353 599
rect -173 565 -161 599
rect 19 565 31 599
rect 211 565 223 599
rect -365 559 -307 565
rect -173 559 -115 565
rect 19 559 77 565
rect 211 559 269 565
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect -365 -565 -307 -559
rect -173 -565 -115 -559
rect 19 -565 77 -559
rect 211 -565 269 -559
rect -365 -599 -353 -565
rect -173 -599 -161 -565
rect 19 -599 31 -565
rect 211 -599 223 -565
rect -365 -605 -307 -599
rect -173 -605 -115 -599
rect 19 -605 77 -599
rect 211 -605 269 -599
<< nwell >>
rect -551 -737 551 737
<< pmos >>
rect -351 118 -321 518
rect -255 118 -225 518
rect -159 118 -129 518
rect -63 118 -33 518
rect 33 118 63 518
rect 129 118 159 518
rect 225 118 255 518
rect 321 118 351 518
rect -351 -518 -321 -118
rect -255 -518 -225 -118
rect -159 -518 -129 -118
rect -63 -518 -33 -118
rect 33 -518 63 -118
rect 129 -518 159 -118
rect 225 -518 255 -118
rect 321 -518 351 -118
<< pdiff >>
rect -413 506 -351 518
rect -413 130 -401 506
rect -367 130 -351 506
rect -413 118 -351 130
rect -321 506 -255 518
rect -321 130 -305 506
rect -271 130 -255 506
rect -321 118 -255 130
rect -225 506 -159 518
rect -225 130 -209 506
rect -175 130 -159 506
rect -225 118 -159 130
rect -129 506 -63 518
rect -129 130 -113 506
rect -79 130 -63 506
rect -129 118 -63 130
rect -33 506 33 518
rect -33 130 -17 506
rect 17 130 33 506
rect -33 118 33 130
rect 63 506 129 518
rect 63 130 79 506
rect 113 130 129 506
rect 63 118 129 130
rect 159 506 225 518
rect 159 130 175 506
rect 209 130 225 506
rect 159 118 225 130
rect 255 506 321 518
rect 255 130 271 506
rect 305 130 321 506
rect 255 118 321 130
rect 351 506 413 518
rect 351 130 367 506
rect 401 130 413 506
rect 351 118 413 130
rect -413 -130 -351 -118
rect -413 -506 -401 -130
rect -367 -506 -351 -130
rect -413 -518 -351 -506
rect -321 -130 -255 -118
rect -321 -506 -305 -130
rect -271 -506 -255 -130
rect -321 -518 -255 -506
rect -225 -130 -159 -118
rect -225 -506 -209 -130
rect -175 -506 -159 -130
rect -225 -518 -159 -506
rect -129 -130 -63 -118
rect -129 -506 -113 -130
rect -79 -506 -63 -130
rect -129 -518 -63 -506
rect -33 -130 33 -118
rect -33 -506 -17 -130
rect 17 -506 33 -130
rect -33 -518 33 -506
rect 63 -130 129 -118
rect 63 -506 79 -130
rect 113 -506 129 -130
rect 63 -518 129 -506
rect 159 -130 225 -118
rect 159 -506 175 -130
rect 209 -506 225 -130
rect 159 -518 225 -506
rect 255 -130 321 -118
rect 255 -506 271 -130
rect 305 -506 321 -130
rect 255 -518 321 -506
rect 351 -130 413 -118
rect 351 -506 367 -130
rect 401 -506 413 -130
rect 351 -518 413 -506
<< pdiffc >>
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
<< nsubdiff >>
rect -515 667 -419 701
rect 419 667 515 701
rect -515 605 -481 667
rect 481 605 515 667
rect -515 -667 -481 -605
rect 481 -667 515 -605
rect -515 -701 -419 -667
rect 419 -701 515 -667
<< nsubdiffcont >>
rect -419 667 419 701
rect -515 -605 -481 605
rect 481 -605 515 605
rect -419 -701 419 -667
<< poly >>
rect -369 599 -303 615
rect -369 565 -353 599
rect -319 565 -303 599
rect -369 549 -303 565
rect -177 599 -111 615
rect -177 565 -161 599
rect -127 565 -111 599
rect -177 549 -111 565
rect 15 599 81 615
rect 15 565 31 599
rect 65 565 81 599
rect 15 549 81 565
rect 207 599 273 615
rect 207 565 223 599
rect 257 565 273 599
rect 207 549 273 565
rect -351 518 -321 549
rect -255 518 -225 544
rect -159 518 -129 549
rect -63 518 -33 544
rect 33 518 63 549
rect 129 518 159 544
rect 225 518 255 549
rect 321 518 351 544
rect -351 92 -321 118
rect -255 87 -225 118
rect -159 92 -129 118
rect -63 87 -33 118
rect 33 92 63 118
rect 129 87 159 118
rect 225 92 255 118
rect 321 87 351 118
rect -273 71 -207 87
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 303 -87 369 -71
rect -351 -118 -321 -92
rect -255 -118 -225 -87
rect -159 -118 -129 -92
rect -63 -118 -33 -87
rect 33 -118 63 -92
rect 129 -118 159 -87
rect 225 -118 255 -92
rect 321 -118 351 -87
rect -351 -549 -321 -518
rect -255 -544 -225 -518
rect -159 -549 -129 -518
rect -63 -544 -33 -518
rect 33 -549 63 -518
rect 129 -544 159 -518
rect 225 -549 255 -518
rect 321 -544 351 -518
rect -369 -565 -303 -549
rect -369 -599 -353 -565
rect -319 -599 -303 -565
rect -369 -615 -303 -599
rect -177 -565 -111 -549
rect -177 -599 -161 -565
rect -127 -599 -111 -565
rect -177 -615 -111 -599
rect 15 -565 81 -549
rect 15 -599 31 -565
rect 65 -599 81 -565
rect 15 -615 81 -599
rect 207 -565 273 -549
rect 207 -599 223 -565
rect 257 -599 273 -565
rect 207 -615 273 -599
<< polycont >>
rect -353 565 -319 599
rect -161 565 -127 599
rect 31 565 65 599
rect 223 565 257 599
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect -353 -599 -319 -565
rect -161 -599 -127 -565
rect 31 -599 65 -565
rect 223 -599 257 -565
<< locali >>
rect -515 667 -419 701
rect 419 667 515 701
rect -515 605 -481 667
rect 481 605 515 667
rect -369 565 -353 599
rect -319 565 -303 599
rect -177 565 -161 599
rect -127 565 -111 599
rect 15 565 31 599
rect 65 565 81 599
rect 207 565 223 599
rect 257 565 273 599
rect -401 506 -367 522
rect -401 114 -367 130
rect -305 506 -271 522
rect -305 114 -271 130
rect -209 506 -175 522
rect -209 114 -175 130
rect -113 506 -79 522
rect -113 114 -79 130
rect -17 506 17 522
rect -17 114 17 130
rect 79 506 113 522
rect 79 114 113 130
rect 175 506 209 522
rect 175 114 209 130
rect 271 506 305 522
rect 271 114 305 130
rect 367 506 401 522
rect 367 114 401 130
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect -401 -130 -367 -114
rect -401 -522 -367 -506
rect -305 -130 -271 -114
rect -305 -522 -271 -506
rect -209 -130 -175 -114
rect -209 -522 -175 -506
rect -113 -130 -79 -114
rect -113 -522 -79 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 79 -130 113 -114
rect 79 -522 113 -506
rect 175 -130 209 -114
rect 175 -522 209 -506
rect 271 -130 305 -114
rect 271 -522 305 -506
rect 367 -130 401 -114
rect 367 -522 401 -506
rect -369 -599 -353 -565
rect -319 -599 -303 -565
rect -177 -599 -161 -565
rect -127 -599 -111 -565
rect 15 -599 31 -565
rect 65 -599 81 -565
rect 207 -599 223 -565
rect 257 -599 273 -565
rect -515 -667 -481 -605
rect 481 -667 515 -605
rect -515 -701 -419 -667
rect 419 -701 515 -667
<< viali >>
rect -353 565 -319 599
rect -161 565 -127 599
rect 31 565 65 599
rect 223 565 257 599
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect -353 -599 -319 -565
rect -161 -599 -127 -565
rect 31 -599 65 -565
rect 223 -599 257 -565
<< metal1 >>
rect -365 599 -307 605
rect -365 565 -353 599
rect -319 565 -307 599
rect -365 559 -307 565
rect -173 599 -115 605
rect -173 565 -161 599
rect -127 565 -115 599
rect -173 559 -115 565
rect 19 599 77 605
rect 19 565 31 599
rect 65 565 77 599
rect 19 559 77 565
rect 211 599 269 605
rect 211 565 223 599
rect 257 565 269 599
rect 211 559 269 565
rect -407 506 -361 518
rect -407 130 -401 506
rect -367 130 -361 506
rect -407 118 -361 130
rect -311 506 -265 518
rect -311 130 -305 506
rect -271 130 -265 506
rect -311 118 -265 130
rect -215 506 -169 518
rect -215 130 -209 506
rect -175 130 -169 506
rect -215 118 -169 130
rect -119 506 -73 518
rect -119 130 -113 506
rect -79 130 -73 506
rect -119 118 -73 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 73 506 119 518
rect 73 130 79 506
rect 113 130 119 506
rect 73 118 119 130
rect 169 506 215 518
rect 169 130 175 506
rect 209 130 215 506
rect 169 118 215 130
rect 265 506 311 518
rect 265 130 271 506
rect 305 130 311 506
rect 265 118 311 130
rect 361 506 407 518
rect 361 130 367 506
rect 401 130 407 506
rect 361 118 407 130
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect -407 -130 -361 -118
rect -407 -506 -401 -130
rect -367 -506 -361 -130
rect -407 -518 -361 -506
rect -311 -130 -265 -118
rect -311 -506 -305 -130
rect -271 -506 -265 -130
rect -311 -518 -265 -506
rect -215 -130 -169 -118
rect -215 -506 -209 -130
rect -175 -506 -169 -130
rect -215 -518 -169 -506
rect -119 -130 -73 -118
rect -119 -506 -113 -130
rect -79 -506 -73 -130
rect -119 -518 -73 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 73 -130 119 -118
rect 73 -506 79 -130
rect 113 -506 119 -130
rect 73 -518 119 -506
rect 169 -130 215 -118
rect 169 -506 175 -130
rect 209 -506 215 -130
rect 169 -518 215 -506
rect 265 -130 311 -118
rect 265 -506 271 -130
rect 305 -506 311 -130
rect 265 -518 311 -506
rect 361 -130 407 -118
rect 361 -506 367 -130
rect 401 -506 407 -130
rect 361 -518 407 -506
rect -365 -565 -307 -559
rect -365 -599 -353 -565
rect -319 -599 -307 -565
rect -365 -605 -307 -599
rect -173 -565 -115 -559
rect -173 -599 -161 -565
rect -127 -599 -115 -565
rect -173 -605 -115 -599
rect 19 -565 77 -559
rect 19 -599 31 -565
rect 65 -599 77 -565
rect 19 -605 77 -599
rect 211 -565 269 -559
rect 211 -599 223 -565
rect 257 -599 269 -565
rect 211 -605 269 -599
<< properties >>
string FIXED_BBOX -498 -684 498 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 2 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
