magic
tech sky130A
magscale 1 2
timestamp 1645179809
<< nwell >>
rect -425 -2691 425 2691
<< pmos >>
rect -229 1672 -29 2472
rect 29 1672 229 2472
rect -229 636 -29 1436
rect 29 636 229 1436
rect -229 -400 -29 400
rect 29 -400 229 400
rect -229 -1436 -29 -636
rect 29 -1436 229 -636
rect -229 -2472 -29 -1672
rect 29 -2472 229 -1672
<< pdiff >>
rect -287 2460 -229 2472
rect -287 1684 -275 2460
rect -241 1684 -229 2460
rect -287 1672 -229 1684
rect -29 2460 29 2472
rect -29 1684 -17 2460
rect 17 1684 29 2460
rect -29 1672 29 1684
rect 229 2460 287 2472
rect 229 1684 241 2460
rect 275 1684 287 2460
rect 229 1672 287 1684
rect -287 1424 -229 1436
rect -287 648 -275 1424
rect -241 648 -229 1424
rect -287 636 -229 648
rect -29 1424 29 1436
rect -29 648 -17 1424
rect 17 648 29 1424
rect -29 636 29 648
rect 229 1424 287 1436
rect 229 648 241 1424
rect 275 648 287 1424
rect 229 636 287 648
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
rect -287 -648 -229 -636
rect -287 -1424 -275 -648
rect -241 -1424 -229 -648
rect -287 -1436 -229 -1424
rect -29 -648 29 -636
rect -29 -1424 -17 -648
rect 17 -1424 29 -648
rect -29 -1436 29 -1424
rect 229 -648 287 -636
rect 229 -1424 241 -648
rect 275 -1424 287 -648
rect 229 -1436 287 -1424
rect -287 -1684 -229 -1672
rect -287 -2460 -275 -1684
rect -241 -2460 -229 -1684
rect -287 -2472 -229 -2460
rect -29 -1684 29 -1672
rect -29 -2460 -17 -1684
rect 17 -2460 29 -1684
rect -29 -2472 29 -2460
rect 229 -1684 287 -1672
rect 229 -2460 241 -1684
rect 275 -2460 287 -1684
rect 229 -2472 287 -2460
<< pdiffc >>
rect -275 1684 -241 2460
rect -17 1684 17 2460
rect 241 1684 275 2460
rect -275 648 -241 1424
rect -17 648 17 1424
rect 241 648 275 1424
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect -275 -1424 -241 -648
rect -17 -1424 17 -648
rect 241 -1424 275 -648
rect -275 -2460 -241 -1684
rect -17 -2460 17 -1684
rect 241 -2460 275 -1684
<< nsubdiff >>
rect -389 2621 -293 2655
rect 293 2621 389 2655
rect -389 2559 -355 2621
rect 355 2559 389 2621
rect -389 -2621 -355 -2559
rect 355 -2621 389 -2559
rect -389 -2655 -293 -2621
rect 293 -2655 389 -2621
<< nsubdiffcont >>
rect -293 2621 293 2655
rect -389 -2559 -355 2559
rect 355 -2559 389 2559
rect -293 -2655 293 -2621
<< poly >>
rect -229 2553 -29 2569
rect -229 2519 -213 2553
rect -45 2519 -29 2553
rect -229 2472 -29 2519
rect 29 2553 229 2569
rect 29 2519 45 2553
rect 213 2519 229 2553
rect 29 2472 229 2519
rect -229 1625 -29 1672
rect -229 1591 -213 1625
rect -45 1591 -29 1625
rect -229 1575 -29 1591
rect 29 1625 229 1672
rect 29 1591 45 1625
rect 213 1591 229 1625
rect 29 1575 229 1591
rect -229 1517 -29 1533
rect -229 1483 -213 1517
rect -45 1483 -29 1517
rect -229 1436 -29 1483
rect 29 1517 229 1533
rect 29 1483 45 1517
rect 213 1483 229 1517
rect 29 1436 229 1483
rect -229 589 -29 636
rect -229 555 -213 589
rect -45 555 -29 589
rect -229 539 -29 555
rect 29 589 229 636
rect 29 555 45 589
rect 213 555 229 589
rect 29 539 229 555
rect -229 481 -29 497
rect -229 447 -213 481
rect -45 447 -29 481
rect -229 400 -29 447
rect 29 481 229 497
rect 29 447 45 481
rect 213 447 229 481
rect 29 400 229 447
rect -229 -447 -29 -400
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect -229 -497 -29 -481
rect 29 -447 229 -400
rect 29 -481 45 -447
rect 213 -481 229 -447
rect 29 -497 229 -481
rect -229 -555 -29 -539
rect -229 -589 -213 -555
rect -45 -589 -29 -555
rect -229 -636 -29 -589
rect 29 -555 229 -539
rect 29 -589 45 -555
rect 213 -589 229 -555
rect 29 -636 229 -589
rect -229 -1483 -29 -1436
rect -229 -1517 -213 -1483
rect -45 -1517 -29 -1483
rect -229 -1533 -29 -1517
rect 29 -1483 229 -1436
rect 29 -1517 45 -1483
rect 213 -1517 229 -1483
rect 29 -1533 229 -1517
rect -229 -1591 -29 -1575
rect -229 -1625 -213 -1591
rect -45 -1625 -29 -1591
rect -229 -1672 -29 -1625
rect 29 -1591 229 -1575
rect 29 -1625 45 -1591
rect 213 -1625 229 -1591
rect 29 -1672 229 -1625
rect -229 -2519 -29 -2472
rect -229 -2553 -213 -2519
rect -45 -2553 -29 -2519
rect -229 -2569 -29 -2553
rect 29 -2519 229 -2472
rect 29 -2553 45 -2519
rect 213 -2553 229 -2519
rect 29 -2569 229 -2553
<< polycont >>
rect -213 2519 -45 2553
rect 45 2519 213 2553
rect -213 1591 -45 1625
rect 45 1591 213 1625
rect -213 1483 -45 1517
rect 45 1483 213 1517
rect -213 555 -45 589
rect 45 555 213 589
rect -213 447 -45 481
rect 45 447 213 481
rect -213 -481 -45 -447
rect 45 -481 213 -447
rect -213 -589 -45 -555
rect 45 -589 213 -555
rect -213 -1517 -45 -1483
rect 45 -1517 213 -1483
rect -213 -1625 -45 -1591
rect 45 -1625 213 -1591
rect -213 -2553 -45 -2519
rect 45 -2553 213 -2519
<< locali >>
rect -389 2621 -293 2655
rect 293 2621 389 2655
rect -389 2559 -355 2621
rect 355 2559 389 2621
rect -229 2519 -213 2553
rect -45 2519 -29 2553
rect 29 2519 45 2553
rect 213 2519 229 2553
rect -275 2460 -241 2476
rect -275 1668 -241 1684
rect -17 2460 17 2476
rect -17 1668 17 1684
rect 241 2460 275 2476
rect 241 1668 275 1684
rect -229 1591 -213 1625
rect -45 1591 -29 1625
rect 29 1591 45 1625
rect 213 1591 229 1625
rect -229 1483 -213 1517
rect -45 1483 -29 1517
rect 29 1483 45 1517
rect 213 1483 229 1517
rect -275 1424 -241 1440
rect -275 632 -241 648
rect -17 1424 17 1440
rect -17 632 17 648
rect 241 1424 275 1440
rect 241 632 275 648
rect -229 555 -213 589
rect -45 555 -29 589
rect 29 555 45 589
rect 213 555 229 589
rect -229 447 -213 481
rect -45 447 -29 481
rect 29 447 45 481
rect 213 447 229 481
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 213 -481 229 -447
rect -229 -589 -213 -555
rect -45 -589 -29 -555
rect 29 -589 45 -555
rect 213 -589 229 -555
rect -275 -648 -241 -632
rect -275 -1440 -241 -1424
rect -17 -648 17 -632
rect -17 -1440 17 -1424
rect 241 -648 275 -632
rect 241 -1440 275 -1424
rect -229 -1517 -213 -1483
rect -45 -1517 -29 -1483
rect 29 -1517 45 -1483
rect 213 -1517 229 -1483
rect -229 -1625 -213 -1591
rect -45 -1625 -29 -1591
rect 29 -1625 45 -1591
rect 213 -1625 229 -1591
rect -275 -1684 -241 -1668
rect -275 -2476 -241 -2460
rect -17 -1684 17 -1668
rect -17 -2476 17 -2460
rect 241 -1684 275 -1668
rect 241 -2476 275 -2460
rect -229 -2553 -213 -2519
rect -45 -2553 -29 -2519
rect 29 -2553 45 -2519
rect 213 -2553 229 -2519
rect -389 -2621 -355 -2559
rect 355 -2621 389 -2559
rect -389 -2655 -293 -2621
rect 293 -2655 389 -2621
<< viali >>
rect -213 2519 -45 2553
rect 45 2519 213 2553
rect -275 1684 -241 2460
rect -17 1684 17 2460
rect 241 1684 275 2460
rect -213 1591 -45 1625
rect 45 1591 213 1625
rect -213 1483 -45 1517
rect 45 1483 213 1517
rect -275 648 -241 1424
rect -17 648 17 1424
rect 241 648 275 1424
rect -213 555 -45 589
rect 45 555 213 589
rect -213 447 -45 481
rect 45 447 213 481
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect -213 -481 -45 -447
rect 45 -481 213 -447
rect -213 -589 -45 -555
rect 45 -589 213 -555
rect -275 -1424 -241 -648
rect -17 -1424 17 -648
rect 241 -1424 275 -648
rect -213 -1517 -45 -1483
rect 45 -1517 213 -1483
rect -213 -1625 -45 -1591
rect 45 -1625 213 -1591
rect -275 -2460 -241 -1684
rect -17 -2460 17 -1684
rect 241 -2460 275 -1684
rect -213 -2553 -45 -2519
rect 45 -2553 213 -2519
<< metal1 >>
rect -225 2553 -33 2559
rect -225 2519 -213 2553
rect -45 2519 -33 2553
rect -225 2513 -33 2519
rect 33 2553 225 2559
rect 33 2519 45 2553
rect 213 2519 225 2553
rect 33 2513 225 2519
rect -281 2460 -235 2472
rect -281 1684 -275 2460
rect -241 1684 -235 2460
rect -281 1672 -235 1684
rect -23 2460 23 2472
rect -23 1684 -17 2460
rect 17 1684 23 2460
rect -23 1672 23 1684
rect 235 2460 281 2472
rect 235 1684 241 2460
rect 275 1684 281 2460
rect 235 1672 281 1684
rect -225 1625 -33 1631
rect -225 1591 -213 1625
rect -45 1591 -33 1625
rect -225 1585 -33 1591
rect 33 1625 225 1631
rect 33 1591 45 1625
rect 213 1591 225 1625
rect 33 1585 225 1591
rect -225 1517 -33 1523
rect -225 1483 -213 1517
rect -45 1483 -33 1517
rect -225 1477 -33 1483
rect 33 1517 225 1523
rect 33 1483 45 1517
rect 213 1483 225 1517
rect 33 1477 225 1483
rect -281 1424 -235 1436
rect -281 648 -275 1424
rect -241 648 -235 1424
rect -281 636 -235 648
rect -23 1424 23 1436
rect -23 648 -17 1424
rect 17 648 23 1424
rect -23 636 23 648
rect 235 1424 281 1436
rect 235 648 241 1424
rect 275 648 281 1424
rect 235 636 281 648
rect -225 589 -33 595
rect -225 555 -213 589
rect -45 555 -33 589
rect -225 549 -33 555
rect 33 589 225 595
rect 33 555 45 589
rect 213 555 225 589
rect 33 549 225 555
rect -225 481 -33 487
rect -225 447 -213 481
rect -45 447 -33 481
rect -225 441 -33 447
rect 33 481 225 487
rect 33 447 45 481
rect 213 447 225 481
rect 33 441 225 447
rect -281 388 -235 400
rect -281 -388 -275 388
rect -241 -388 -235 388
rect -281 -400 -235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 235 388 281 400
rect 235 -388 241 388
rect 275 -388 281 388
rect 235 -400 281 -388
rect -225 -447 -33 -441
rect -225 -481 -213 -447
rect -45 -481 -33 -447
rect -225 -487 -33 -481
rect 33 -447 225 -441
rect 33 -481 45 -447
rect 213 -481 225 -447
rect 33 -487 225 -481
rect -225 -555 -33 -549
rect -225 -589 -213 -555
rect -45 -589 -33 -555
rect -225 -595 -33 -589
rect 33 -555 225 -549
rect 33 -589 45 -555
rect 213 -589 225 -555
rect 33 -595 225 -589
rect -281 -648 -235 -636
rect -281 -1424 -275 -648
rect -241 -1424 -235 -648
rect -281 -1436 -235 -1424
rect -23 -648 23 -636
rect -23 -1424 -17 -648
rect 17 -1424 23 -648
rect -23 -1436 23 -1424
rect 235 -648 281 -636
rect 235 -1424 241 -648
rect 275 -1424 281 -648
rect 235 -1436 281 -1424
rect -225 -1483 -33 -1477
rect -225 -1517 -213 -1483
rect -45 -1517 -33 -1483
rect -225 -1523 -33 -1517
rect 33 -1483 225 -1477
rect 33 -1517 45 -1483
rect 213 -1517 225 -1483
rect 33 -1523 225 -1517
rect -225 -1591 -33 -1585
rect -225 -1625 -213 -1591
rect -45 -1625 -33 -1591
rect -225 -1631 -33 -1625
rect 33 -1591 225 -1585
rect 33 -1625 45 -1591
rect 213 -1625 225 -1591
rect 33 -1631 225 -1625
rect -281 -1684 -235 -1672
rect -281 -2460 -275 -1684
rect -241 -2460 -235 -1684
rect -281 -2472 -235 -2460
rect -23 -1684 23 -1672
rect -23 -2460 -17 -1684
rect 17 -2460 23 -1684
rect -23 -2472 23 -2460
rect 235 -1684 281 -1672
rect 235 -2460 241 -1684
rect 275 -2460 281 -1684
rect 235 -2472 281 -2460
rect -225 -2519 -33 -2513
rect -225 -2553 -213 -2519
rect -45 -2553 -33 -2519
rect -225 -2559 -33 -2553
rect 33 -2519 225 -2513
rect 33 -2553 45 -2519
rect 213 -2553 225 -2519
rect 33 -2559 225 -2553
<< properties >>
string FIXED_BBOX -372 -2638 372 2638
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 1 m 5 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
