magic
tech sky130A
magscale 1 2
timestamp 1645531774
<< nwell >>
rect -4473 -591 -3807 591
rect -3553 -591 -2887 591
rect -2633 -591 -1967 591
rect -1713 -591 -1047 591
rect -793 -591 -127 591
rect 127 -591 793 591
rect 1047 -591 1713 591
rect 1967 -591 2633 591
rect 2887 -591 3553 591
rect 3807 -591 4473 591
<< pwell >>
rect -4583 591 4583 701
rect -4583 -591 -4473 591
rect -3807 -591 -3553 591
rect -2887 -591 -2633 591
rect -1967 -591 -1713 591
rect -1047 -591 -793 591
rect -127 -591 127 591
rect 793 -591 1047 591
rect 1713 -591 1967 591
rect 2633 -591 2887 591
rect 3553 -591 3807 591
rect 4473 -591 4583 591
rect -4583 -701 4583 -591
<< varactor >>
rect -4340 -500 -3940 500
rect -3420 -500 -3020 500
rect -2500 -500 -2100 500
rect -1580 -500 -1180 500
rect -660 -500 -260 500
rect 260 -500 660 500
rect 1180 -500 1580 500
rect 2100 -500 2500 500
rect 3020 -500 3420 500
rect 3940 -500 4340 500
<< psubdiff >>
rect -4547 631 -4451 665
rect 4451 631 4547 665
rect -4547 569 -4513 631
rect 4513 569 4547 631
rect -4547 -631 -4513 -569
rect 4513 -631 4547 -569
rect -4547 -665 -4451 -631
rect 4451 -665 4547 -631
<< nsubdiff >>
rect -4437 476 -4340 500
rect -4437 -476 -4425 476
rect -4391 -476 -4340 476
rect -4437 -500 -4340 -476
rect -3940 476 -3843 500
rect -3940 -476 -3889 476
rect -3855 -476 -3843 476
rect -3940 -500 -3843 -476
rect -3517 476 -3420 500
rect -3517 -476 -3505 476
rect -3471 -476 -3420 476
rect -3517 -500 -3420 -476
rect -3020 476 -2923 500
rect -3020 -476 -2969 476
rect -2935 -476 -2923 476
rect -3020 -500 -2923 -476
rect -2597 476 -2500 500
rect -2597 -476 -2585 476
rect -2551 -476 -2500 476
rect -2597 -500 -2500 -476
rect -2100 476 -2003 500
rect -2100 -476 -2049 476
rect -2015 -476 -2003 476
rect -2100 -500 -2003 -476
rect -1677 476 -1580 500
rect -1677 -476 -1665 476
rect -1631 -476 -1580 476
rect -1677 -500 -1580 -476
rect -1180 476 -1083 500
rect -1180 -476 -1129 476
rect -1095 -476 -1083 476
rect -1180 -500 -1083 -476
rect -757 476 -660 500
rect -757 -476 -745 476
rect -711 -476 -660 476
rect -757 -500 -660 -476
rect -260 476 -163 500
rect -260 -476 -209 476
rect -175 -476 -163 476
rect -260 -500 -163 -476
rect 163 476 260 500
rect 163 -476 175 476
rect 209 -476 260 476
rect 163 -500 260 -476
rect 660 476 757 500
rect 660 -476 711 476
rect 745 -476 757 476
rect 660 -500 757 -476
rect 1083 476 1180 500
rect 1083 -476 1095 476
rect 1129 -476 1180 476
rect 1083 -500 1180 -476
rect 1580 476 1677 500
rect 1580 -476 1631 476
rect 1665 -476 1677 476
rect 1580 -500 1677 -476
rect 2003 476 2100 500
rect 2003 -476 2015 476
rect 2049 -476 2100 476
rect 2003 -500 2100 -476
rect 2500 476 2597 500
rect 2500 -476 2551 476
rect 2585 -476 2597 476
rect 2500 -500 2597 -476
rect 2923 476 3020 500
rect 2923 -476 2935 476
rect 2969 -476 3020 476
rect 2923 -500 3020 -476
rect 3420 476 3517 500
rect 3420 -476 3471 476
rect 3505 -476 3517 476
rect 3420 -500 3517 -476
rect 3843 476 3940 500
rect 3843 -476 3855 476
rect 3889 -476 3940 476
rect 3843 -500 3940 -476
rect 4340 476 4437 500
rect 4340 -476 4391 476
rect 4425 -476 4437 476
rect 4340 -500 4437 -476
<< psubdiffcont >>
rect -4451 631 4451 665
rect -4547 -569 -4513 569
rect 4513 -569 4547 569
rect -4451 -665 4451 -631
<< nsubdiffcont >>
rect -4425 -476 -4391 476
rect -3889 -476 -3855 476
rect -3505 -476 -3471 476
rect -2969 -476 -2935 476
rect -2585 -476 -2551 476
rect -2049 -476 -2015 476
rect -1665 -476 -1631 476
rect -1129 -476 -1095 476
rect -745 -476 -711 476
rect -209 -476 -175 476
rect 175 -476 209 476
rect 711 -476 745 476
rect 1095 -476 1129 476
rect 1631 -476 1665 476
rect 2015 -476 2049 476
rect 2551 -476 2585 476
rect 2935 -476 2969 476
rect 3471 -476 3505 476
rect 3855 -476 3889 476
rect 4391 -476 4425 476
<< poly >>
rect -4340 572 -3940 588
rect -4340 538 -4324 572
rect -3956 538 -3940 572
rect -4340 500 -3940 538
rect -3420 572 -3020 588
rect -3420 538 -3404 572
rect -3036 538 -3020 572
rect -3420 500 -3020 538
rect -2500 572 -2100 588
rect -2500 538 -2484 572
rect -2116 538 -2100 572
rect -2500 500 -2100 538
rect -1580 572 -1180 588
rect -1580 538 -1564 572
rect -1196 538 -1180 572
rect -1580 500 -1180 538
rect -660 572 -260 588
rect -660 538 -644 572
rect -276 538 -260 572
rect -660 500 -260 538
rect 260 572 660 588
rect 260 538 276 572
rect 644 538 660 572
rect 260 500 660 538
rect 1180 572 1580 588
rect 1180 538 1196 572
rect 1564 538 1580 572
rect 1180 500 1580 538
rect 2100 572 2500 588
rect 2100 538 2116 572
rect 2484 538 2500 572
rect 2100 500 2500 538
rect 3020 572 3420 588
rect 3020 538 3036 572
rect 3404 538 3420 572
rect 3020 500 3420 538
rect 3940 572 4340 588
rect 3940 538 3956 572
rect 4324 538 4340 572
rect 3940 500 4340 538
rect -4340 -538 -3940 -500
rect -4340 -572 -4324 -538
rect -3956 -572 -3940 -538
rect -4340 -588 -3940 -572
rect -3420 -538 -3020 -500
rect -3420 -572 -3404 -538
rect -3036 -572 -3020 -538
rect -3420 -588 -3020 -572
rect -2500 -538 -2100 -500
rect -2500 -572 -2484 -538
rect -2116 -572 -2100 -538
rect -2500 -588 -2100 -572
rect -1580 -538 -1180 -500
rect -1580 -572 -1564 -538
rect -1196 -572 -1180 -538
rect -1580 -588 -1180 -572
rect -660 -538 -260 -500
rect -660 -572 -644 -538
rect -276 -572 -260 -538
rect -660 -588 -260 -572
rect 260 -538 660 -500
rect 260 -572 276 -538
rect 644 -572 660 -538
rect 260 -588 660 -572
rect 1180 -538 1580 -500
rect 1180 -572 1196 -538
rect 1564 -572 1580 -538
rect 1180 -588 1580 -572
rect 2100 -538 2500 -500
rect 2100 -572 2116 -538
rect 2484 -572 2500 -538
rect 2100 -588 2500 -572
rect 3020 -538 3420 -500
rect 3020 -572 3036 -538
rect 3404 -572 3420 -538
rect 3020 -588 3420 -572
rect 3940 -538 4340 -500
rect 3940 -572 3956 -538
rect 4324 -572 4340 -538
rect 3940 -588 4340 -572
<< polycont >>
rect -4324 538 -3956 572
rect -3404 538 -3036 572
rect -2484 538 -2116 572
rect -1564 538 -1196 572
rect -644 538 -276 572
rect 276 538 644 572
rect 1196 538 1564 572
rect 2116 538 2484 572
rect 3036 538 3404 572
rect 3956 538 4324 572
rect -4324 -572 -3956 -538
rect -3404 -572 -3036 -538
rect -2484 -572 -2116 -538
rect -1564 -572 -1196 -538
rect -644 -572 -276 -538
rect 276 -572 644 -538
rect 1196 -572 1564 -538
rect 2116 -572 2484 -538
rect 3036 -572 3404 -538
rect 3956 -572 4324 -538
<< locali >>
rect -4547 631 -4451 665
rect 4451 631 4547 665
rect -4547 569 -4513 631
rect -4340 538 -4324 572
rect -3956 538 -3940 572
rect -3420 538 -3404 572
rect -3036 538 -3020 572
rect -2500 538 -2484 572
rect -2116 538 -2100 572
rect -1580 538 -1564 572
rect -1196 538 -1180 572
rect -660 538 -644 572
rect -276 538 -260 572
rect 260 538 276 572
rect 644 538 660 572
rect 1180 538 1196 572
rect 1564 538 1580 572
rect 2100 538 2116 572
rect 2484 538 2500 572
rect 3020 538 3036 572
rect 3404 538 3420 572
rect 3940 538 3956 572
rect 4324 538 4340 572
rect 4513 569 4547 631
rect -4425 476 -4391 492
rect -4425 -492 -4391 -476
rect -3889 476 -3855 492
rect -3889 -492 -3855 -476
rect -3505 476 -3471 492
rect -3505 -492 -3471 -476
rect -2969 476 -2935 492
rect -2969 -492 -2935 -476
rect -2585 476 -2551 492
rect -2585 -492 -2551 -476
rect -2049 476 -2015 492
rect -2049 -492 -2015 -476
rect -1665 476 -1631 492
rect -1665 -492 -1631 -476
rect -1129 476 -1095 492
rect -1129 -492 -1095 -476
rect -745 476 -711 492
rect -745 -492 -711 -476
rect -209 476 -175 492
rect -209 -492 -175 -476
rect 175 476 209 492
rect 175 -492 209 -476
rect 711 476 745 492
rect 711 -492 745 -476
rect 1095 476 1129 492
rect 1095 -492 1129 -476
rect 1631 476 1665 492
rect 1631 -492 1665 -476
rect 2015 476 2049 492
rect 2015 -492 2049 -476
rect 2551 476 2585 492
rect 2551 -492 2585 -476
rect 2935 476 2969 492
rect 2935 -492 2969 -476
rect 3471 476 3505 492
rect 3471 -492 3505 -476
rect 3855 476 3889 492
rect 3855 -492 3889 -476
rect 4391 476 4425 492
rect 4391 -492 4425 -476
rect -4547 -631 -4513 -569
rect -4340 -572 -4324 -538
rect -3956 -572 -3940 -538
rect -3420 -572 -3404 -538
rect -3036 -572 -3020 -538
rect -2500 -572 -2484 -538
rect -2116 -572 -2100 -538
rect -1580 -572 -1564 -538
rect -1196 -572 -1180 -538
rect -660 -572 -644 -538
rect -276 -572 -260 -538
rect 260 -572 276 -538
rect 644 -572 660 -538
rect 1180 -572 1196 -538
rect 1564 -572 1580 -538
rect 2100 -572 2116 -538
rect 2484 -572 2500 -538
rect 3020 -572 3036 -538
rect 3404 -572 3420 -538
rect 3940 -572 3956 -538
rect 4324 -572 4340 -538
rect 4513 -631 4547 -569
rect -4547 -665 -4451 -631
rect 4451 -665 4547 -631
<< viali >>
rect -4324 538 -3956 572
rect -3404 538 -3036 572
rect -2484 538 -2116 572
rect -1564 538 -1196 572
rect -644 538 -276 572
rect 276 538 644 572
rect 1196 538 1564 572
rect 2116 538 2484 572
rect 3036 538 3404 572
rect 3956 538 4324 572
rect -4425 -476 -4391 476
rect -3889 -476 -3855 476
rect -3505 -476 -3471 476
rect -2969 -476 -2935 476
rect -2585 -476 -2551 476
rect -2049 -476 -2015 476
rect -1665 -476 -1631 476
rect -1129 -476 -1095 476
rect -745 -476 -711 476
rect -209 -476 -175 476
rect 175 -476 209 476
rect 711 -476 745 476
rect 1095 -476 1129 476
rect 1631 -476 1665 476
rect 2015 -476 2049 476
rect 2551 -476 2585 476
rect 2935 -476 2969 476
rect 3471 -476 3505 476
rect 3855 -476 3889 476
rect 4391 -476 4425 476
rect -4324 -572 -3956 -538
rect -3404 -572 -3036 -538
rect -2484 -572 -2116 -538
rect -1564 -572 -1196 -538
rect -644 -572 -276 -538
rect 276 -572 644 -538
rect 1196 -572 1564 -538
rect 2116 -572 2484 -538
rect 3036 -572 3404 -538
rect 3956 -572 4324 -538
<< metal1 >>
rect -4336 572 -3944 578
rect -4336 538 -4324 572
rect -3956 538 -3944 572
rect -4336 532 -3944 538
rect -3416 572 -3024 578
rect -3416 538 -3404 572
rect -3036 538 -3024 572
rect -3416 532 -3024 538
rect -2496 572 -2104 578
rect -2496 538 -2484 572
rect -2116 538 -2104 572
rect -2496 532 -2104 538
rect -1576 572 -1184 578
rect -1576 538 -1564 572
rect -1196 538 -1184 572
rect -1576 532 -1184 538
rect -656 572 -264 578
rect -656 538 -644 572
rect -276 538 -264 572
rect -656 532 -264 538
rect 264 572 656 578
rect 264 538 276 572
rect 644 538 656 572
rect 264 532 656 538
rect 1184 572 1576 578
rect 1184 538 1196 572
rect 1564 538 1576 572
rect 1184 532 1576 538
rect 2104 572 2496 578
rect 2104 538 2116 572
rect 2484 538 2496 572
rect 2104 532 2496 538
rect 3024 572 3416 578
rect 3024 538 3036 572
rect 3404 538 3416 572
rect 3024 532 3416 538
rect 3944 572 4336 578
rect 3944 538 3956 572
rect 4324 538 4336 572
rect 3944 532 4336 538
rect -4431 476 -4385 488
rect -4431 -476 -4425 476
rect -4391 -476 -4385 476
rect -4431 -488 -4385 -476
rect -3895 476 -3849 488
rect -3895 -476 -3889 476
rect -3855 -476 -3849 476
rect -3895 -488 -3849 -476
rect -3511 476 -3465 488
rect -3511 -476 -3505 476
rect -3471 -476 -3465 476
rect -3511 -488 -3465 -476
rect -2975 476 -2929 488
rect -2975 -476 -2969 476
rect -2935 -476 -2929 476
rect -2975 -488 -2929 -476
rect -2591 476 -2545 488
rect -2591 -476 -2585 476
rect -2551 -476 -2545 476
rect -2591 -488 -2545 -476
rect -2055 476 -2009 488
rect -2055 -476 -2049 476
rect -2015 -476 -2009 476
rect -2055 -488 -2009 -476
rect -1671 476 -1625 488
rect -1671 -476 -1665 476
rect -1631 -476 -1625 476
rect -1671 -488 -1625 -476
rect -1135 476 -1089 488
rect -1135 -476 -1129 476
rect -1095 -476 -1089 476
rect -1135 -488 -1089 -476
rect -751 476 -705 488
rect -751 -476 -745 476
rect -711 -476 -705 476
rect -751 -488 -705 -476
rect -215 476 -169 488
rect -215 -476 -209 476
rect -175 -476 -169 476
rect -215 -488 -169 -476
rect 169 476 215 488
rect 169 -476 175 476
rect 209 -476 215 476
rect 169 -488 215 -476
rect 705 476 751 488
rect 705 -476 711 476
rect 745 -476 751 476
rect 705 -488 751 -476
rect 1089 476 1135 488
rect 1089 -476 1095 476
rect 1129 -476 1135 476
rect 1089 -488 1135 -476
rect 1625 476 1671 488
rect 1625 -476 1631 476
rect 1665 -476 1671 476
rect 1625 -488 1671 -476
rect 2009 476 2055 488
rect 2009 -476 2015 476
rect 2049 -476 2055 476
rect 2009 -488 2055 -476
rect 2545 476 2591 488
rect 2545 -476 2551 476
rect 2585 -476 2591 476
rect 2545 -488 2591 -476
rect 2929 476 2975 488
rect 2929 -476 2935 476
rect 2969 -476 2975 476
rect 2929 -488 2975 -476
rect 3465 476 3511 488
rect 3465 -476 3471 476
rect 3505 -476 3511 476
rect 3465 -488 3511 -476
rect 3849 476 3895 488
rect 3849 -476 3855 476
rect 3889 -476 3895 476
rect 3849 -488 3895 -476
rect 4385 476 4431 488
rect 4385 -476 4391 476
rect 4425 -476 4431 476
rect 4385 -488 4431 -476
rect -4336 -538 -3944 -532
rect -4336 -572 -4324 -538
rect -3956 -572 -3944 -538
rect -4336 -578 -3944 -572
rect -3416 -538 -3024 -532
rect -3416 -572 -3404 -538
rect -3036 -572 -3024 -538
rect -3416 -578 -3024 -572
rect -2496 -538 -2104 -532
rect -2496 -572 -2484 -538
rect -2116 -572 -2104 -538
rect -2496 -578 -2104 -572
rect -1576 -538 -1184 -532
rect -1576 -572 -1564 -538
rect -1196 -572 -1184 -538
rect -1576 -578 -1184 -572
rect -656 -538 -264 -532
rect -656 -572 -644 -538
rect -276 -572 -264 -538
rect -656 -578 -264 -572
rect 264 -538 656 -532
rect 264 -572 276 -538
rect 644 -572 656 -538
rect 264 -578 656 -572
rect 1184 -538 1576 -532
rect 1184 -572 1196 -538
rect 1564 -572 1576 -538
rect 1184 -578 1576 -572
rect 2104 -538 2496 -532
rect 2104 -572 2116 -538
rect 2484 -572 2496 -538
rect 2104 -578 2496 -572
rect 3024 -538 3416 -532
rect 3024 -572 3036 -538
rect 3404 -572 3416 -538
rect 3024 -578 3416 -572
rect 3944 -538 4336 -532
rect 3944 -572 3956 -538
rect 4324 -572 4336 -538
rect 3944 -578 4336 -572
<< properties >>
string FIXED_BBOX -4530 -648 4530 648
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 5 l 2 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
