magic
tech sky130B
magscale 1 2
timestamp 1653928699
<< nwell >>
rect -1290 4230 -1060 4450
<< pwell >>
rect 4450 1180 4770 1210
rect 4960 1180 7980 1210
rect 4460 670 4780 700
rect 4960 670 7970 700
rect 8670 -450 8860 -400
rect 8380 -500 8910 -480
rect 8380 -660 9150 -500
<< locali >>
rect 1420 1400 1520 2140
rect 850 1310 2090 1400
rect 1430 560 1510 1310
rect -640 -960 -530 -890
rect -630 -1600 -510 -1530
rect -110 -1590 -30 -1520
<< viali >>
rect -30 -1670 40 -1490
<< metal1 >>
rect -8730 6580 -8410 6630
rect -6060 6590 -5660 6620
rect -6210 6380 -6200 6540
rect -6140 6380 -6130 6540
rect -6020 6380 -6010 6540
rect -5950 6380 -5940 6540
rect -5830 6380 -5820 6540
rect -5760 6380 -5750 6540
rect -6120 6140 -6110 6300
rect -6050 6140 -6040 6300
rect -5930 6140 -5920 6300
rect -5860 6140 -5850 6300
rect -9040 5760 -8980 6080
rect -8700 6050 -8380 6100
rect -5690 6090 -5660 6590
rect -4170 6580 -3860 6630
rect -2820 6580 -2510 6630
rect 5210 6580 5610 6630
rect 6540 6580 6940 6630
rect 8430 6590 8820 6620
rect 8280 6380 8290 6540
rect 8350 6380 8360 6540
rect 8470 6380 8480 6540
rect 8540 6380 8550 6540
rect 8660 6380 8670 6540
rect 8730 6380 8740 6540
rect 8370 6140 8380 6300
rect 8440 6140 8450 6300
rect 8560 6140 8570 6300
rect 8630 6140 8640 6300
rect -7950 5760 -7890 6080
rect -6860 5760 -6800 6080
rect -6150 6060 -5280 6090
rect -8740 4940 -8460 4990
rect -7620 4940 -7340 4990
rect -6550 4940 -6270 4990
rect -9040 4120 -8980 4440
rect -8740 4410 -8420 4460
rect -7950 4120 -7890 4440
rect -7650 4410 -7330 4460
rect -6860 4120 -6800 4440
rect -6550 4410 -6270 4460
rect -6130 4370 -6120 4450
rect -5850 4370 -5840 4450
rect -5770 4120 -5710 4440
rect -8710 3300 -8430 3350
rect -7620 3300 -7300 3350
rect -6540 3300 -6260 3350
rect -6170 3300 -5420 3350
rect -8700 2770 -8420 2820
rect -7620 2770 -7300 2820
rect -6530 2770 -6250 2820
rect -6170 2770 -5850 2820
rect -5320 2550 -5280 6060
rect -5000 5770 -4950 6070
rect -4140 6050 -3830 6100
rect -3660 5770 -3610 6070
rect -2790 6050 -2480 6100
rect -2320 5790 -2270 6090
rect 4140 6050 7980 6100
rect 8790 6090 8820 6590
rect 10120 6580 10450 6630
rect 11200 6580 11530 6630
rect 8080 6060 8820 6090
rect 4380 5730 4430 6050
rect 5720 5730 5770 6050
rect 7060 5730 7110 6050
rect -4150 4940 -3860 4990
rect -2790 4940 -2500 4990
rect 5210 4940 5610 4990
rect 6550 4940 6950 4990
rect -5000 4150 -4950 4450
rect -4160 4410 -3870 4460
rect -3660 4140 -3610 4440
rect -2810 4410 -2520 4460
rect -2320 4140 -2270 4440
rect 4140 4410 7980 4460
rect 4380 4090 4430 4410
rect 5720 4090 5770 4410
rect 7060 4090 7110 4410
rect -4160 3300 -3870 3350
rect -2890 3300 -2480 3350
rect -1520 3300 -1110 3350
rect -120 3300 180 3350
rect 2550 3300 2850 3350
rect 3850 3300 4150 3350
rect 5250 3300 5550 3350
rect 6600 3300 6900 3350
rect -4100 2770 -3810 2820
rect -2860 2770 -2450 2820
rect -1510 2770 -1100 2820
rect -110 2770 190 2820
rect 970 2730 980 2800
rect 1180 2730 1190 2800
rect 1750 2720 1760 2820
rect 1970 2720 1980 2820
rect 2590 2770 2890 2820
rect 3850 2770 7610 2820
rect 8080 2550 8120 6060
rect 9810 5770 9870 6070
rect 10130 6050 10460 6100
rect 10900 5780 10960 6080
rect 11230 6050 11560 6100
rect 11990 5780 12050 6080
rect 8350 5220 8380 5280
rect 10120 4940 10450 4990
rect 11230 4940 11560 4990
rect 8160 4500 8170 4660
rect 8240 4500 8250 4660
rect 8720 4120 8780 4440
rect 9810 4150 9870 4450
rect 10120 4410 10450 4460
rect 10900 4150 10960 4450
rect 11220 4410 11550 4460
rect 11990 4150 12050 4450
rect 9040 3300 9370 3350
rect 10140 3300 10470 3350
rect 11190 3300 11520 3350
rect 9030 2770 9360 2820
rect 10140 2770 10470 2820
rect 11220 2770 11550 2820
rect -5320 2510 -800 2550
rect -810 2470 -800 2510
rect -720 2510 8120 2550
rect -720 2470 -710 2510
rect 8810 2400 8820 2440
rect -6320 2370 8820 2400
rect 8900 2370 8910 2440
rect -9530 1180 -6650 1210
rect -6320 1180 -6290 2370
rect -6000 2290 9030 2320
rect -9530 670 -6650 700
rect -9270 -400 -9240 -80
rect -8570 -400 -8540 -70
rect -7870 -400 -7840 -70
rect -9530 -430 -7280 -400
rect -7170 -410 -7140 -70
rect -6000 -410 -5970 2290
rect 2910 2210 2920 2250
rect -1270 2180 2920 2210
rect 2990 2180 3000 2250
rect -1270 1880 -1190 2180
rect -160 2140 4160 2150
rect -170 2070 -160 2140
rect -90 2120 4160 2140
rect -90 2070 -80 2120
rect 1020 1990 1440 2060
rect -1280 1810 -1270 1880
rect -1190 1810 -1180 1880
rect 1110 1790 1120 1960
rect 1190 1790 1200 1960
rect -5490 1580 200 1660
rect -5490 1180 -5400 1580
rect -1280 1370 -1270 1440
rect -1190 1370 -1180 1440
rect -170 1370 -160 1440
rect -90 1370 -80 1440
rect -5100 1180 -1580 1210
rect -1270 1180 -1190 1370
rect -830 1270 -820 1370
rect -730 1270 -720 1370
rect -5100 670 -1570 700
rect -4880 -410 -4850 -20
rect -4180 -410 -4150 -20
rect -6390 -440 -6120 -410
rect -6000 -440 -5810 -410
rect -5090 -440 -3650 -410
rect -3480 -440 -3450 -20
rect -9530 -940 -7280 -910
rect -6390 -920 -6350 -440
rect -6220 -640 -6210 -480
rect -6150 -640 -6140 -480
rect -5900 -640 -5890 -480
rect -5830 -640 -5820 -480
rect -6310 -880 -6300 -720
rect -6240 -880 -6230 -720
rect -6120 -880 -6110 -720
rect -6050 -880 -6040 -720
rect -6390 -950 -6220 -920
rect -5090 -950 -3650 -920
rect -6260 -1120 -6220 -950
rect -820 -960 -790 1270
rect -400 1190 -390 1250
rect -240 1190 -230 1250
rect -160 1180 -90 1370
rect 120 1220 200 1580
rect 950 1560 960 1730
rect 1030 1560 1040 1730
rect 1270 1560 1280 1730
rect 1350 1560 1360 1730
rect 1390 1530 1440 1990
rect 1020 1460 1440 1530
rect 1510 1990 1930 2060
rect 4100 1990 4160 2120
rect 1510 1530 1560 1990
rect 1750 1790 1760 1960
rect 1830 1790 1840 1960
rect 4090 1930 4100 1990
rect 4160 1930 4170 1990
rect 8820 1960 8830 2020
rect 8890 1960 8900 2020
rect 1590 1560 1600 1730
rect 1670 1560 1680 1730
rect 1910 1560 1920 1730
rect 1990 1560 2000 1730
rect 1510 1460 1930 1530
rect 2620 1400 8280 1440
rect 2620 1220 2720 1400
rect 2910 1300 2920 1360
rect 2990 1300 3000 1360
rect 120 1180 2720 1220
rect 2920 1180 2990 1300
rect 3120 1240 3130 1320
rect 3280 1240 3290 1320
rect 4090 1310 4100 1370
rect 4160 1310 4170 1370
rect 3040 1180 3090 1220
rect 3120 1200 3290 1240
rect 4100 1180 4160 1310
rect 4450 1180 4770 1210
rect 4960 1180 7980 1210
rect 8210 1180 8280 1400
rect 4460 670 4780 700
rect 4960 670 7970 700
rect 410 -430 440 -80
rect 570 -440 840 -410
rect 1110 -420 1140 -80
rect 1370 -440 1400 -410
rect 1390 -470 1400 -440
rect 1560 -470 1570 -410
rect 1810 -430 1840 -80
rect 1980 -440 2250 -410
rect 2510 -430 2540 -80
rect 6400 -410 6430 -40
rect 7100 -410 7130 -40
rect 6150 -440 7720 -410
rect 7800 -440 7830 -40
rect 8440 -420 8450 -360
rect 8570 -420 8580 -360
rect 8840 -400 8880 1960
rect 9000 1200 9030 2290
rect 9000 1180 9090 1200
rect 9390 1180 11890 1210
rect 9390 670 11890 700
rect 8670 -450 8880 -400
rect 9990 -410 10020 -80
rect 10690 -410 10720 -80
rect 11390 -410 11420 -80
rect 12090 -410 12120 -80
rect 9140 -450 9330 -420
rect 9760 -440 12260 -410
rect 9080 -660 9090 -490
rect 9150 -660 9160 -490
rect -720 -770 -430 -720
rect -820 -990 -730 -960
rect -650 -980 -640 -840
rect -580 -980 -570 -840
rect -6280 -1200 -6270 -1120
rect -6190 -1200 -6180 -1120
rect -820 -1460 -790 -990
rect -470 -1050 -430 -770
rect 8990 -890 9000 -720
rect 9060 -890 9070 -720
rect 9180 -890 9190 -720
rect 9250 -890 9260 -720
rect 560 -950 830 -920
rect 1290 -950 1560 -920
rect 1980 -950 2250 -920
rect 6180 -950 7750 -920
rect 9290 -930 9330 -450
rect -720 -1100 -430 -1050
rect -470 -1180 -430 -1100
rect 9050 -960 9330 -930
rect 9750 -950 12230 -920
rect -470 -1230 -130 -1180
rect 9050 -1230 9090 -960
rect -470 -1380 -420 -1230
rect -700 -1430 -420 -1380
rect -250 -1430 -240 -1260
rect -180 -1430 -170 -1260
rect 9020 -1350 9030 -1230
rect 9140 -1350 9150 -1230
rect -820 -1500 -710 -1460
rect -710 -1640 -700 -1590
rect -640 -1650 -630 -1510
rect -570 -1650 -560 -1510
rect -470 -1690 -420 -1430
rect -36 -1490 46 -1478
rect -340 -1660 -330 -1490
rect -270 -1660 -260 -1490
rect -150 -1660 -140 -1490
rect -80 -1660 -70 -1490
rect -36 -1670 -30 -1490
rect 40 -1670 46 -1490
rect -36 -1682 46 -1670
rect -710 -1710 -220 -1690
rect -960 -1740 -220 -1710
rect -1030 -1870 -1020 -1800
rect -960 -1870 -930 -1740
rect -280 -1760 -220 -1740
rect 20 -1760 30 -1740
rect -280 -1800 30 -1760
rect 20 -1830 30 -1800
rect 110 -1830 120 -1740
<< via1 >>
rect -6200 6380 -6140 6540
rect -6010 6380 -5950 6540
rect -5820 6380 -5760 6540
rect -6110 6140 -6050 6300
rect -5920 6140 -5860 6300
rect 8290 6380 8350 6540
rect 8480 6380 8540 6540
rect 8670 6380 8730 6540
rect 8380 6140 8440 6300
rect 8570 6140 8630 6300
rect -6120 4370 -5850 4450
rect 980 2730 1180 2800
rect 1760 2720 1970 2820
rect 8170 4500 8240 4660
rect -800 2470 -720 2550
rect 8820 2370 8900 2440
rect 2920 2180 2990 2250
rect -160 2070 -90 2140
rect -1270 1810 -1190 1880
rect 1120 1790 1190 1960
rect -1270 1370 -1190 1440
rect -160 1370 -90 1440
rect -820 1270 -730 1370
rect -6210 -640 -6150 -480
rect -5890 -640 -5830 -480
rect -6300 -880 -6240 -720
rect -6110 -880 -6050 -720
rect -390 1190 -240 1250
rect 960 1560 1030 1730
rect 1280 1560 1350 1730
rect 1760 1790 1830 1960
rect 4100 1930 4160 1990
rect 8830 1960 8890 2020
rect 1600 1560 1670 1730
rect 1920 1560 1990 1730
rect 2920 1300 2990 1360
rect 3130 1240 3280 1320
rect 4100 1310 4160 1370
rect 1400 -470 1560 -410
rect 8450 -420 8570 -360
rect 9090 -660 9150 -490
rect -640 -980 -580 -840
rect -6270 -1200 -6190 -1120
rect 9000 -890 9060 -720
rect 9190 -890 9250 -720
rect -240 -1430 -180 -1260
rect 9030 -1350 9140 -1230
rect -630 -1650 -570 -1510
rect -330 -1660 -270 -1490
rect -140 -1660 -80 -1490
rect -1020 -1870 -960 -1800
rect 30 -1830 110 -1740
<< metal2 >>
rect -6280 7560 -5770 7570
rect -9460 7200 -6280 7560
rect -6310 7190 -6280 7200
rect -5770 7530 -570 7560
rect 8470 7550 9100 7560
rect -5770 7190 -1200 7530
rect -5770 7040 -5220 7190
rect -1200 7050 -570 7060
rect -6280 7030 -5220 7040
rect -6240 6778 -5220 7030
rect -5790 6550 -5220 6778
rect -6200 6540 -5220 6550
rect -1990 6540 -1800 6550
rect -9350 6520 -6590 6540
rect -9350 6380 -8000 6520
rect -7920 6380 -6590 6520
rect -6140 6380 -6010 6540
rect -5950 6380 -5820 6540
rect -5760 6380 -5220 6540
rect -5120 6530 -1990 6540
rect -5120 6390 -5110 6530
rect -8000 6370 -7920 6380
rect -6200 6370 -6140 6380
rect -6010 6370 -5950 6380
rect -5820 6370 -5220 6380
rect -4920 6390 -1990 6530
rect -1800 6390 -1350 6540
rect -1990 6380 -1800 6390
rect -5110 6370 -4920 6380
rect -6120 6300 -5850 6310
rect -9350 6290 -6590 6300
rect -9350 6140 -7780 6290
rect -7200 6140 -6590 6290
rect -7780 6130 -7200 6140
rect -6120 6120 -5850 6130
rect -5790 5920 -5220 6370
rect -4800 6300 -4610 6310
rect -1660 6300 -1470 6310
rect -4990 6150 -4800 6300
rect -4610 6150 -1660 6300
rect -4800 6140 -4610 6150
rect -1660 6140 -1470 6150
rect -1030 5920 -570 7050
rect -9450 5560 -570 5920
rect -6240 5550 -6170 5560
rect -5760 5550 -570 5560
rect -9350 4890 -6590 4900
rect -5110 4890 -4920 4900
rect -1990 4890 -1800 4900
rect -9350 4750 -8000 4890
rect -7920 4750 -6590 4890
rect -9350 4740 -6590 4750
rect -5120 4740 -5110 4890
rect -4920 4740 -1990 4890
rect -1800 4740 -1600 4890
rect -5110 4730 -4920 4740
rect -1990 4730 -1800 4740
rect -6120 4660 -5850 4670
rect -9350 4650 -6590 4660
rect -9350 4500 -7780 4650
rect -7200 4500 -6590 4650
rect -5800 4660 -4610 4670
rect -1660 4660 -1470 4670
rect -5800 4510 -4800 4660
rect -4610 4510 -1660 4660
rect -5800 4500 -4610 4510
rect -1660 4500 -1470 4510
rect -7780 4490 -7200 4500
rect -6120 4450 -5850 4500
rect -6120 4360 -5850 4370
rect -1030 4290 -570 5550
rect 2990 7540 3620 7550
rect 3620 7180 8470 7540
rect 2990 7060 3620 7070
rect 9100 7190 11940 7550
rect 2990 5910 3450 7060
rect 8470 6550 9100 7080
rect 4260 6540 4450 6550
rect 8290 6540 9100 6550
rect 4450 6530 8020 6540
rect 4450 6390 7390 6530
rect 4260 6380 4450 6390
rect 7580 6390 8020 6530
rect 7390 6370 7580 6380
rect 8350 6380 8480 6540
rect 8540 6380 8670 6540
rect 8730 6380 9100 6540
rect 9380 6540 9540 6550
rect 8290 6370 9100 6380
rect 9370 6370 9380 6530
rect 11770 6530 11960 6540
rect 9540 6380 11770 6530
rect 9540 6370 11960 6380
rect 7700 6300 7890 6310
rect 4590 6290 4780 6300
rect 5970 6290 6190 6300
rect 4380 6140 4590 6290
rect 4780 6140 5970 6290
rect 6190 6150 7700 6290
rect 8380 6300 8630 6310
rect 7890 6150 7900 6290
rect 6190 6140 7900 6150
rect 8440 6140 8570 6150
rect 4590 6130 4780 6140
rect 5970 6130 6190 6140
rect 8380 6130 8630 6140
rect 8680 5910 9100 6370
rect 9380 6360 9540 6370
rect 9670 6310 9830 6320
rect 9460 6140 9670 6300
rect 12110 6300 12300 6310
rect 9830 6290 12020 6300
rect 9830 6150 10660 6290
rect 11050 6150 12020 6290
rect 9830 6140 12020 6150
rect 12110 6140 12300 6150
rect 9670 6130 9830 6140
rect 2990 5880 11920 5910
rect 2990 5590 6420 5880
rect 6990 5590 8700 5880
rect 2990 5580 8700 5590
rect 2990 5550 8320 5580
rect 9300 5710 11920 5880
rect 9300 5570 11930 5710
rect 8700 5550 11930 5570
rect -5290 4280 -240 4290
rect 2990 4280 3450 5550
rect 4260 4900 4450 4910
rect 9380 4900 9540 4910
rect 4450 4890 8030 4900
rect 4450 4750 7390 4890
rect 4260 4740 4450 4750
rect 7580 4750 8030 4890
rect 7390 4730 7580 4740
rect 9370 4730 9380 4890
rect 11770 4890 11960 4900
rect 9540 4740 11770 4890
rect 9540 4730 11960 4740
rect 9380 4720 9540 4730
rect 9670 4670 9830 4680
rect 7700 4660 7890 4670
rect 8170 4660 8240 4670
rect 4590 4650 4780 4660
rect 5970 4650 6190 4660
rect 7200 4650 7700 4660
rect 4380 4500 4590 4650
rect 4780 4500 5970 4650
rect 6190 4510 7700 4650
rect 7890 4510 8170 4660
rect 6190 4500 8170 4510
rect 8240 4650 8690 4660
rect 8240 4510 8390 4650
rect 8590 4510 8690 4650
rect 9460 4510 9670 4670
rect 8240 4500 8690 4510
rect 9830 4660 12020 4670
rect 9830 4520 10660 4660
rect 11050 4520 12020 4660
rect 9830 4510 12020 4520
rect 12110 4660 12300 4670
rect 12110 4500 12300 4510
rect 4590 4490 4780 4500
rect 5970 4490 6190 4500
rect 8170 4490 8240 4500
rect 9670 4490 9830 4500
rect -9470 4270 8120 4280
rect -9470 3940 -5710 4270
rect -5280 4260 8120 4270
rect 9200 4260 11900 4270
rect -5280 4240 11900 4260
rect -5280 4080 8700 4240
rect -5280 3940 -600 4080
rect -9470 3920 -600 3940
rect -5730 3910 -600 3920
rect -480 3910 6420 4080
rect 6990 3930 8700 4080
rect 9300 4080 11900 4240
rect 9300 3930 11940 4080
rect 6990 3910 8150 3930
rect 8700 3920 11940 3930
rect 8780 3910 11940 3920
rect -600 3900 -480 3910
rect 6420 3900 6990 3910
rect -1990 3260 -1800 3270
rect 4260 3260 4450 3270
rect 9380 3260 9540 3270
rect -5110 3250 -1990 3260
rect -9340 3240 -6590 3250
rect -9340 3100 -8000 3240
rect -7920 3100 -6590 3240
rect -9340 3090 -6590 3100
rect -4920 3110 -1990 3250
rect -1800 3110 -1590 3260
rect 4450 3250 8020 3260
rect 4450 3110 7390 3250
rect -1990 3100 -1800 3110
rect 4260 3100 4450 3110
rect 7580 3110 8020 3250
rect -5110 3090 -4920 3100
rect 7390 3090 7580 3100
rect 9540 3250 12220 3260
rect 9540 3100 11770 3250
rect 11960 3100 12220 3250
rect 9540 3090 12220 3100
rect 9380 3080 9540 3090
rect 9670 3030 9830 3040
rect -5700 3020 -5460 3030
rect -4800 3020 -4610 3030
rect -1660 3020 -1470 3030
rect -9340 3010 -6590 3020
rect -9340 2860 -7780 3010
rect -7200 2860 -6590 3010
rect -7780 2850 -7200 2860
rect -5700 2850 -5460 2860
rect -5000 2870 -4800 3020
rect -4610 2870 -1660 3020
rect 1190 3020 1320 3030
rect 7700 3020 7890 3030
rect -5000 2860 -4610 2870
rect -1660 2860 -1470 2870
rect -9380 1220 -6330 1230
rect -9380 990 -7780 1220
rect -7200 990 -6330 1220
rect -9380 980 -6330 990
rect -5700 1140 -5450 1150
rect -5000 1140 -4780 2860
rect -800 2550 -720 2560
rect -1270 1880 -1190 1890
rect -1270 1440 -1190 1810
rect -800 1410 -720 2470
rect -1270 1360 -1190 1370
rect -820 1370 -720 1410
rect -820 1260 -730 1270
rect -390 1250 -240 3000
rect 980 2800 1190 3010
rect 1180 2730 1190 2800
rect 980 2640 1190 2730
rect 1530 3010 1860 3020
rect 4590 3010 4780 3020
rect 5970 3010 6190 3020
rect 7650 3010 7700 3020
rect 1860 2860 1970 2920
rect 3130 2890 3280 3010
rect 1530 2850 1970 2860
rect 980 2630 1320 2640
rect 1760 2820 1970 2850
rect 3100 2820 3280 2890
rect 4390 2860 4590 3010
rect 4780 2860 5970 3010
rect 6190 2870 7700 3010
rect 8390 3020 8590 3030
rect 7890 2870 7910 3010
rect 6190 2860 7910 2870
rect 9460 2860 9670 3030
rect 9830 3020 12300 3030
rect 9830 2860 10660 3020
rect 11050 2870 12110 3020
rect 11050 2860 12300 2870
rect 4590 2850 4780 2860
rect 5970 2850 6190 2860
rect 7650 2850 7870 2860
rect 8390 2850 8590 2860
rect -160 2140 -90 2150
rect -160 1440 -90 2070
rect 980 1960 1190 2630
rect 980 1790 1120 1960
rect 1120 1780 1190 1790
rect 1760 1960 1970 2720
rect 1830 1790 1970 1960
rect 1760 1780 1970 1790
rect 2920 2250 2990 2260
rect 960 1730 1030 1740
rect 1280 1730 1350 1740
rect 1600 1730 1670 1740
rect 1920 1730 1990 1740
rect 1030 1560 1280 1730
rect 1350 1560 1600 1730
rect 1670 1560 1920 1730
rect 960 1550 1990 1560
rect -160 1360 -90 1370
rect -390 1140 -240 1190
rect 1360 1140 1580 1550
rect 2920 1360 2990 2180
rect 2920 1290 2990 1300
rect 3130 1320 3280 2820
rect 9470 2540 12300 2860
rect 8820 2440 8900 2450
rect 8820 2360 8900 2370
rect 8840 2030 8880 2360
rect 8830 2020 8890 2030
rect 4100 1990 4160 2000
rect 8830 1950 8890 1960
rect 4100 1370 4160 1930
rect 11750 1340 12300 2540
rect 4100 1300 4160 1310
rect -5700 1130 -1260 1140
rect -5700 990 -5000 1130
rect -4860 990 -3660 1130
rect -3520 990 -1260 1130
rect -5700 980 -1260 990
rect -410 980 -170 1140
rect 300 980 2640 1140
rect 3130 1020 3280 1240
rect 9180 1150 12300 1340
rect 5970 1140 6190 1150
rect 6810 1140 7220 1150
rect 9180 1140 10840 1150
rect 3320 1130 3340 1140
rect 4190 980 5970 1140
rect 6190 1130 8460 1140
rect 6190 990 6270 1130
rect 6410 990 7660 1130
rect 7880 990 8460 1130
rect 6190 980 8460 990
rect 9170 1130 10840 1140
rect 9170 990 9870 1130
rect 10010 990 10840 1130
rect 11230 1130 12300 1150
rect 11230 990 11870 1130
rect 12010 1050 12300 1130
rect 12010 990 12200 1050
rect 9170 980 12200 990
rect 5970 970 6190 980
rect 6810 970 7220 980
rect -9490 890 -6270 900
rect -9490 750 -8200 890
rect -8110 750 -6270 890
rect -9490 740 -6270 750
rect -5090 890 -1190 900
rect -5090 750 -4790 890
rect -4650 750 -3390 890
rect -3250 750 -1190 890
rect -5090 740 -1190 750
rect 250 740 2560 900
rect 4080 890 8040 900
rect 4080 750 6510 890
rect 6650 750 7890 890
rect 8030 750 8040 890
rect 4080 740 8040 750
rect 9090 890 12010 900
rect 9090 750 10130 890
rect 10270 750 12010 890
rect 9090 740 12010 750
rect 12160 890 12300 900
rect 12160 740 12300 750
rect -990 100 3030 120
rect 3180 100 5470 120
rect 5720 100 9000 120
rect -9130 90 9000 100
rect -9130 -70 12310 90
rect -9130 -240 12320 -70
rect -9130 -290 -930 -240
rect -7780 -390 -7200 -380
rect -9390 -620 -7780 -390
rect -7200 -620 -7030 -390
rect -9390 -630 -7030 -620
rect -6860 -410 -6330 -290
rect -9260 -720 -6960 -710
rect -9260 -860 -8200 -720
rect -8110 -860 -6960 -720
rect -9260 -870 -6960 -860
rect -6860 -1000 -6850 -410
rect -6350 -710 -6330 -410
rect -3050 -420 -930 -290
rect -6210 -480 -6150 -470
rect -5890 -480 -5830 -470
rect -6150 -640 -5890 -480
rect -5830 -490 -5450 -480
rect -5830 -640 -5700 -490
rect -5000 -490 -3340 -480
rect -4860 -630 -3660 -490
rect -3520 -630 -3340 -490
rect -5000 -640 -3340 -630
rect -6210 -650 -6150 -640
rect -5890 -650 -5830 -640
rect -5700 -650 -5450 -640
rect -6350 -720 -6050 -710
rect -6350 -880 -6300 -720
rect -6240 -880 -6110 -720
rect -5040 -730 -3250 -720
rect -5090 -870 -4790 -730
rect -4650 -870 -3390 -730
rect -5090 -880 -3250 -870
rect -6350 -890 -6050 -880
rect -6350 -1000 -6330 -890
rect -6860 -1510 -6330 -1000
rect -3050 -1000 -3020 -420
rect -2140 -830 -930 -420
rect 1400 -410 1560 -400
rect 1270 -460 1400 -450
rect 2860 -420 3710 -240
rect 1560 -460 1630 -450
rect -600 -540 -480 -530
rect -600 -670 -480 -660
rect -50 -640 310 -480
rect 430 -630 1270 -470
rect 1630 -630 2440 -470
rect 430 -640 2440 -630
rect -600 -830 -510 -670
rect -2140 -1000 -2110 -830
rect -3050 -1030 -2110 -1000
rect -6270 -1120 -6190 -1110
rect -6270 -1210 -6190 -1200
rect -3050 -1510 -2120 -1030
rect -9140 -1900 -2120 -1510
rect -1150 -1490 -930 -830
rect -640 -840 -510 -830
rect -580 -930 -510 -840
rect -50 -870 130 -640
rect -640 -990 -580 -980
rect 200 -880 2330 -720
rect -50 -1250 130 -1230
rect -240 -1260 130 -1250
rect -180 -1430 130 -1260
rect -240 -1440 130 -1430
rect 2860 -990 2900 -420
rect 3680 -990 3710 -420
rect -330 -1490 -270 -1480
rect -140 -1490 -80 -1480
rect -1150 -1510 -330 -1490
rect -1150 -1650 -630 -1510
rect -570 -1650 -330 -1510
rect -1150 -1660 -330 -1650
rect -270 -1660 -140 -1490
rect -80 -1530 200 -1490
rect 2860 -1530 3710 -990
rect -80 -1660 3710 -1530
rect -330 -1670 3710 -1660
rect 30 -1740 110 -1730
rect -1020 -1800 -960 -1790
rect 30 -1840 110 -1830
rect 190 -1860 3710 -1670
rect 5350 -430 6070 -240
rect 9010 -280 9650 -240
rect 5350 -1000 5360 -430
rect 6040 -1000 6070 -430
rect 8450 -360 8570 -350
rect 6890 -480 7220 -470
rect 8450 -480 8570 -420
rect 9290 -420 9650 -280
rect 6270 -490 6890 -480
rect 6410 -630 6890 -490
rect 6270 -640 6890 -630
rect 7220 -490 7940 -480
rect 7220 -630 7660 -490
rect 7800 -630 7940 -490
rect 7220 -640 7940 -630
rect 8380 -490 9150 -480
rect 8380 -630 8390 -490
rect 8590 -630 9090 -490
rect 6890 -650 7220 -640
rect 8380 -660 9090 -630
rect 9090 -670 9150 -660
rect 9290 -710 9310 -420
rect 9000 -720 9310 -710
rect 6180 -730 7850 -720
rect 6180 -870 6510 -730
rect 6650 -870 7850 -730
rect 6180 -880 7850 -870
rect 7890 -730 8030 -720
rect 7890 -880 8030 -870
rect 9060 -890 9190 -720
rect 9250 -890 9310 -720
rect 9000 -900 9310 -890
rect 5350 -1530 6070 -1000
rect 9290 -1000 9310 -900
rect 9630 -1000 9650 -420
rect 9870 -490 12220 -480
rect 10010 -630 10840 -490
rect 11230 -630 11870 -490
rect 12010 -630 12220 -490
rect 9870 -640 12220 -630
rect 9770 -730 12320 -720
rect 9770 -870 10130 -730
rect 10270 -870 12160 -730
rect 12300 -870 12320 -730
rect 9770 -880 12320 -870
rect 9030 -1230 9140 -1220
rect 9030 -1360 9140 -1350
rect 9290 -1530 9650 -1000
rect 5350 -1860 12330 -1530
rect 190 -1870 3440 -1860
rect -1020 -1880 -960 -1870
<< via2 >>
rect -6280 7040 -5770 7560
rect -1200 7060 -570 7530
rect -8000 6380 -7920 6520
rect -5110 6380 -4920 6530
rect -1990 6390 -1800 6540
rect -7780 6140 -7200 6290
rect -6120 6140 -6110 6300
rect -6110 6140 -6050 6300
rect -6050 6140 -5920 6300
rect -5920 6140 -5860 6300
rect -5860 6140 -5850 6300
rect -6120 6130 -5850 6140
rect -4800 6150 -4610 6300
rect -1660 6150 -1470 6300
rect -8000 4750 -7920 4890
rect -5110 4740 -4920 4890
rect -1990 4740 -1800 4890
rect -7780 4500 -7200 4650
rect -6120 4500 -5850 4660
rect -4800 4510 -4610 4660
rect -1660 4510 -1470 4660
rect 2990 7070 3620 7540
rect 8470 7080 9100 7550
rect 4260 6390 4450 6540
rect 7390 6380 7580 6530
rect 9380 6370 9540 6540
rect 11770 6380 11960 6530
rect 4590 6140 4780 6290
rect 5970 6140 6190 6290
rect 7700 6150 7890 6300
rect 8390 6150 8440 6300
rect 8440 6150 8570 6300
rect 8570 6150 8590 6300
rect 9670 6140 9830 6310
rect 10660 6150 11050 6290
rect 12110 6150 12300 6300
rect 6420 5590 6990 5880
rect 8700 5570 9300 5880
rect 4260 4750 4450 4900
rect 7390 4740 7580 4890
rect 9380 4730 9540 4900
rect 11770 4740 11960 4890
rect 4590 4500 4780 4650
rect 5970 4500 6190 4650
rect 7700 4510 7890 4660
rect 8390 4510 8590 4650
rect 9670 4500 9830 4670
rect 10660 4520 11050 4660
rect 12110 4510 12300 4660
rect -5710 3940 -5280 4270
rect -600 3910 -480 4080
rect 6420 3910 6990 4080
rect 8700 3930 9300 4240
rect -8000 3100 -7920 3240
rect -5110 3100 -4920 3250
rect -1990 3110 -1800 3260
rect 4260 3110 4450 3260
rect 7390 3100 7580 3250
rect 9380 3090 9540 3260
rect 11770 3100 11960 3250
rect -7780 2860 -7200 3010
rect -5700 2860 -5460 3020
rect -4800 2870 -4610 3020
rect -1660 2870 -1470 3020
rect -7780 990 -7200 1220
rect 1190 2640 1320 3020
rect 1530 2860 1860 3010
rect 4590 2860 4780 3010
rect 5970 2860 6190 3010
rect 7700 2870 7890 3020
rect 8390 2860 8590 3020
rect 9670 2860 9830 3030
rect 10660 2860 11050 3020
rect 12110 2870 12300 3020
rect -5000 990 -4860 1130
rect -3660 990 -3520 1130
rect 5970 980 6190 1140
rect 6270 990 6410 1130
rect 7660 990 7880 1130
rect 9870 990 10010 1130
rect 10840 990 11230 1150
rect 11870 990 12010 1130
rect -8200 750 -8110 890
rect -4790 750 -4650 890
rect -3390 750 -3250 890
rect 6510 750 6650 890
rect 7890 750 8030 890
rect 10130 750 10270 890
rect 12160 750 12300 890
rect -7780 -620 -7200 -390
rect -8200 -860 -8110 -720
rect -6850 -1000 -6350 -410
rect -5700 -640 -5450 -490
rect -5000 -630 -4860 -490
rect -3660 -630 -3520 -490
rect -4790 -870 -4650 -730
rect -3390 -870 -3250 -730
rect -3020 -1000 -2140 -420
rect 1270 -470 1400 -460
rect 1400 -470 1560 -460
rect 1560 -470 1630 -460
rect -600 -660 -480 -540
rect 1270 -630 1630 -470
rect -6270 -1200 -6190 -1120
rect -50 -1230 130 -870
rect 2900 -990 3680 -420
rect -1020 -1870 -960 -1800
rect 30 -1830 110 -1740
rect 5360 -1000 6040 -430
rect 6270 -630 6410 -490
rect 6890 -640 7220 -480
rect 7660 -630 7800 -490
rect 8390 -630 8590 -490
rect 6510 -870 6650 -730
rect 7890 -870 8030 -730
rect 9310 -1000 9630 -420
rect 9870 -630 10010 -490
rect 10840 -630 11230 -490
rect 11870 -630 12010 -490
rect 10130 -870 10270 -730
rect 12160 -870 12300 -730
rect 9030 -1350 9140 -1230
<< metal3 >>
rect -6290 7560 -5760 7565
rect -6290 7040 -6280 7560
rect -5770 7300 -5360 7560
rect 8460 7550 9110 7555
rect 2980 7540 3630 7545
rect -1210 7530 -560 7535
rect -5770 7040 -5280 7300
rect -1210 7060 -1200 7530
rect -570 7060 -560 7530
rect 2980 7070 2990 7540
rect 3620 7070 3630 7540
rect 8460 7080 8470 7550
rect 9100 7080 9300 7550
rect 8460 7075 9300 7080
rect 2980 7065 3630 7070
rect -1210 7055 -560 7060
rect -6290 6980 -5280 7040
rect -8010 6520 -7910 6525
rect -8010 6380 -8000 6520
rect -7920 6380 -7910 6520
rect -8010 6375 -7910 6380
rect -8000 4895 -7920 6375
rect -6130 6300 -5840 6305
rect -7780 6295 -7200 6300
rect -7790 6290 -7190 6295
rect -7790 6140 -7780 6290
rect -7200 6140 -7190 6290
rect -7790 6135 -7190 6140
rect -8010 4890 -7910 4895
rect -8010 4750 -8000 4890
rect -7920 4750 -7910 4890
rect -8010 4745 -7910 4750
rect -8000 3245 -7920 4745
rect -7780 4655 -7200 6135
rect -6130 6130 -6120 6300
rect -5850 6130 -5840 6300
rect -6130 6125 -5840 6130
rect -6120 4665 -5840 6125
rect -6130 4660 -5840 4665
rect -7790 4650 -7190 4655
rect -7790 4500 -7780 4650
rect -7200 4500 -7190 4650
rect -7790 4495 -7190 4500
rect -6130 4500 -6120 4660
rect -5850 4500 -5840 4660
rect -6130 4495 -5840 4500
rect -8010 3240 -7910 3245
rect -8010 3100 -8000 3240
rect -7920 3100 -7910 3240
rect -8010 3095 -7910 3100
rect -7780 3015 -7200 4495
rect -5710 4275 -5280 6980
rect -2000 6540 -1790 6545
rect -5110 6535 -4920 6540
rect -5120 6530 -4910 6535
rect -5120 6380 -5110 6530
rect -4920 6380 -4910 6530
rect -5120 6375 -4910 6380
rect -2000 6390 -1990 6540
rect -1800 6390 -1790 6540
rect -2000 6385 -1790 6390
rect 4250 6540 4460 6545
rect 4250 6390 4260 6540
rect 4450 6390 4460 6540
rect 7390 6535 7580 6550
rect 4250 6385 4460 6390
rect 7380 6530 7590 6535
rect -5110 4895 -4920 6375
rect -4800 6305 -4610 6310
rect -4810 6300 -4600 6305
rect -4810 6150 -4800 6300
rect -4610 6150 -4600 6300
rect -4810 6145 -4600 6150
rect -5120 4890 -4910 4895
rect -5120 4740 -5110 4890
rect -4920 4740 -4910 4890
rect -5120 4735 -4910 4740
rect -5720 4270 -5270 4275
rect -5720 3940 -5710 4270
rect -5280 3940 -5270 4270
rect -5720 3935 -5270 3940
rect -5110 3255 -4920 4735
rect -4800 4665 -4610 6145
rect -2000 4895 -1810 6385
rect -1670 6300 -1460 6305
rect -1670 6150 -1660 6300
rect -1470 6150 -1460 6300
rect -1670 6145 -1460 6150
rect -2000 4890 -1790 4895
rect -2000 4740 -1990 4890
rect -1800 4740 -1790 4890
rect -2000 4735 -1790 4740
rect -4810 4660 -4600 4665
rect -4810 4510 -4800 4660
rect -4610 4510 -4600 4660
rect -4810 4505 -4600 4510
rect -5120 3250 -4910 3255
rect -5120 3100 -5110 3250
rect -4920 3100 -4910 3250
rect -5120 3095 -4910 3100
rect -5700 3025 -5450 3030
rect -4800 3025 -4610 4505
rect -2000 3265 -1810 4735
rect -1660 4665 -1470 6145
rect 4260 4905 4450 6385
rect 7380 6380 7390 6530
rect 7580 6380 7590 6530
rect 7380 6375 7590 6380
rect 4580 6290 4790 6295
rect 4580 6140 4590 6290
rect 4780 6140 4790 6290
rect 4580 6135 4790 6140
rect 5960 6290 6200 6295
rect 5960 6140 5970 6290
rect 6190 6140 6200 6290
rect 5960 6135 6200 6140
rect 4250 4900 4460 4905
rect 4250 4750 4260 4900
rect 4450 4750 4460 4900
rect 4250 4745 4460 4750
rect -1670 4660 -1460 4665
rect -1670 4510 -1660 4660
rect -1470 4510 -1460 4660
rect -1670 4505 -1460 4510
rect -2000 3260 -1790 3265
rect -2000 3110 -1990 3260
rect -1800 3110 -1790 3260
rect -2000 3105 -1790 3110
rect -1660 3025 -1470 4505
rect -610 4080 -470 4085
rect -610 3910 -600 4080
rect -480 3910 -470 4080
rect -610 3905 -470 3910
rect -5710 3020 -5450 3025
rect -7790 3010 -7190 3015
rect -7790 2860 -7780 3010
rect -7200 2860 -7190 3010
rect -7790 2855 -7190 2860
rect -5710 2860 -5700 3020
rect -5460 2860 -5450 3020
rect -4810 3020 -4600 3025
rect -4810 2870 -4800 3020
rect -4610 2870 -4600 3020
rect -4810 2865 -4600 2870
rect -1670 3020 -1460 3025
rect -1670 2870 -1660 3020
rect -1470 2870 -1460 3020
rect -1670 2865 -1460 2870
rect -5710 2855 -5450 2860
rect -7780 1225 -7200 2855
rect -7790 1220 -7190 1225
rect -7790 990 -7780 1220
rect -7200 990 -7190 1220
rect -7790 985 -7190 990
rect -8200 895 -8110 900
rect -8210 890 -8100 895
rect -8210 750 -8200 890
rect -8110 750 -8100 890
rect -8210 745 -8100 750
rect -8200 -715 -8110 745
rect -7780 -385 -7200 985
rect -7790 -390 -7190 -385
rect -7790 -620 -7780 -390
rect -7200 -620 -7190 -390
rect -7790 -625 -7190 -620
rect -6860 -410 -6340 -405
rect -7780 -630 -7200 -625
rect -8210 -720 -8100 -715
rect -8210 -860 -8200 -720
rect -8110 -860 -8100 -720
rect -8210 -865 -8100 -860
rect -8200 -870 -8110 -865
rect -6860 -1000 -6850 -410
rect -6350 -1000 -6340 -410
rect -5700 -485 -5450 2855
rect -5000 1135 -4860 1140
rect -3660 1135 -3520 1140
rect -5010 1130 -4850 1135
rect -5010 990 -5000 1130
rect -4860 990 -4850 1130
rect -5010 985 -4850 990
rect -3670 1130 -3510 1135
rect -3670 990 -3660 1130
rect -3520 990 -3510 1130
rect -3670 985 -3510 990
rect -5000 -485 -4860 985
rect -4790 895 -4650 900
rect -4800 890 -4640 895
rect -4800 750 -4790 890
rect -4650 750 -4640 890
rect -4800 745 -4640 750
rect -5710 -490 -5440 -485
rect -5710 -640 -5700 -490
rect -5450 -640 -5440 -490
rect -5010 -490 -4850 -485
rect -5010 -630 -5000 -490
rect -4860 -630 -4850 -490
rect -5010 -635 -4850 -630
rect -5000 -640 -4860 -635
rect -5710 -645 -5440 -640
rect -4790 -725 -4650 745
rect -3660 -485 -3520 985
rect -3390 895 -3250 900
rect -3400 890 -3240 895
rect -3400 750 -3390 890
rect -3250 750 -3240 890
rect -3400 745 -3240 750
rect -3670 -490 -3510 -485
rect -3670 -630 -3660 -490
rect -3520 -630 -3510 -490
rect -3670 -635 -3510 -630
rect -3660 -640 -3520 -635
rect -3390 -725 -3250 745
rect -3030 -420 -2130 -415
rect -4800 -730 -4640 -725
rect -4800 -870 -4790 -730
rect -4650 -870 -4640 -730
rect -4800 -875 -4640 -870
rect -3400 -730 -3240 -725
rect -3400 -870 -3390 -730
rect -3250 -870 -3240 -730
rect -3400 -875 -3240 -870
rect -4790 -880 -4650 -875
rect -3390 -880 -3250 -875
rect -6860 -1005 -6340 -1000
rect -3030 -1000 -3020 -420
rect -2140 -1000 -2130 -420
rect -600 -535 -480 3905
rect 4260 3265 4450 4745
rect 4590 4655 4780 6135
rect 5970 4655 6190 6135
rect 6410 5880 7000 5885
rect 6410 5590 6420 5880
rect 6990 5590 7000 5880
rect 6410 5585 7000 5590
rect 4580 4650 4790 4655
rect 4580 4500 4590 4650
rect 4780 4500 4790 4650
rect 4580 4495 4790 4500
rect 5960 4650 6200 4655
rect 5960 4500 5970 4650
rect 6190 4500 6200 4650
rect 5960 4495 6200 4500
rect 4250 3260 4460 3265
rect 4250 3110 4260 3260
rect 4450 3110 4460 3260
rect 4250 3105 4460 3110
rect 1180 3020 1330 3025
rect 1180 2640 1190 3020
rect 1320 2640 1330 3020
rect 1520 2640 1530 3030
rect 1670 3015 1680 3030
rect 4590 3015 4780 4495
rect 5970 3015 6190 4495
rect 6420 4085 6990 5585
rect 7390 4895 7580 6375
rect 7700 6305 7890 6310
rect 7690 6300 7900 6305
rect 7690 6150 7700 6300
rect 7890 6150 7900 6300
rect 7690 6145 7900 6150
rect 8380 6300 8600 6305
rect 8380 6150 8390 6300
rect 8590 6150 8600 6300
rect 8380 6145 8600 6150
rect 7380 4890 7590 4895
rect 7380 4740 7390 4890
rect 7580 4740 7590 4890
rect 7380 4735 7590 4740
rect 6410 4080 7000 4085
rect 6410 3910 6420 4080
rect 6990 3910 7000 4080
rect 6410 3905 7000 3910
rect 1670 3010 1870 3015
rect 1860 2860 1870 3010
rect 1670 2855 1870 2860
rect 4580 3010 4790 3015
rect 4580 2860 4590 3010
rect 4780 2860 4790 3010
rect 4580 2855 4790 2860
rect 5960 3010 6200 3015
rect 5960 2860 5970 3010
rect 6190 2860 6200 3010
rect 5960 2855 6200 2860
rect 1670 2640 1680 2855
rect 1180 2635 1330 2640
rect 5970 1145 6190 2855
rect 6420 2720 6990 3905
rect 7390 3255 7580 4735
rect 7700 4665 7890 6145
rect 7690 4660 7900 4665
rect 7690 4510 7700 4660
rect 7890 4510 7900 4660
rect 8390 4655 8590 6145
rect 8700 5885 9300 7075
rect 9370 6540 9550 6545
rect 9370 6370 9380 6540
rect 9540 6370 9550 6540
rect 11760 6530 11970 6535
rect 11760 6380 11770 6530
rect 11960 6380 11970 6530
rect 11760 6375 11970 6380
rect 9370 6365 9550 6370
rect 8690 5880 9310 5885
rect 8690 5570 8700 5880
rect 9300 5570 9310 5880
rect 8690 5565 9310 5570
rect 7690 4505 7900 4510
rect 8380 4650 8600 4655
rect 8380 4510 8390 4650
rect 8590 4510 8600 4650
rect 8380 4505 8600 4510
rect 7380 3250 7590 3255
rect 7380 3100 7390 3250
rect 7580 3100 7590 3250
rect 7380 3095 7590 3100
rect 7700 3040 7890 4505
rect 8700 4245 9300 5565
rect 9380 4905 9540 6365
rect 9660 6310 9840 6315
rect 9660 6140 9670 6310
rect 9830 6140 9840 6310
rect 10650 6290 11060 6295
rect 10650 6150 10660 6290
rect 11050 6150 11060 6290
rect 10650 6145 11060 6150
rect 9660 6135 9840 6140
rect 9370 4900 9550 4905
rect 9370 4730 9380 4900
rect 9540 4730 9550 4900
rect 9370 4725 9550 4730
rect 8690 4240 9310 4245
rect 8690 3930 8700 4240
rect 9300 3930 9310 4240
rect 8690 3925 9310 3930
rect 9380 3265 9540 4725
rect 9670 4675 9830 6135
rect 9660 4670 9840 4675
rect 9660 4500 9670 4670
rect 9830 4500 9840 4670
rect 10660 4665 11050 6145
rect 11770 4895 11960 6375
rect 12100 6300 12310 6305
rect 12100 6150 12110 6300
rect 12300 6150 12310 6300
rect 12100 6145 12310 6150
rect 11760 4890 11970 4895
rect 11760 4740 11770 4890
rect 11960 4740 11970 4890
rect 11760 4735 11970 4740
rect 10650 4660 11060 4665
rect 10650 4520 10660 4660
rect 11050 4520 11060 4660
rect 10650 4515 11060 4520
rect 9660 4495 9840 4500
rect 9370 3260 9550 3265
rect 9370 3090 9380 3260
rect 9540 3090 9550 3260
rect 9370 3085 9550 3090
rect 7700 3025 7900 3040
rect 9670 3035 9830 4495
rect 9660 3030 9840 3035
rect 8390 3025 8590 3030
rect 7690 3020 7900 3025
rect 7690 2870 7700 3020
rect 7890 2870 7900 3020
rect 7690 2865 7900 2870
rect 5960 1140 6200 1145
rect 7700 1140 7900 2865
rect 8380 3020 8600 3025
rect 8380 2860 8390 3020
rect 8590 2860 8600 3020
rect 8380 2855 8600 2860
rect 9660 2860 9670 3030
rect 9830 2860 9840 3030
rect 10660 3025 11050 4515
rect 11770 3255 11960 4735
rect 12110 4665 12300 6145
rect 12100 4660 12310 4665
rect 12100 4510 12110 4660
rect 12300 4510 12310 4660
rect 12100 4505 12310 4510
rect 11760 3250 11970 3255
rect 11760 3100 11770 3250
rect 11960 3100 11970 3250
rect 11760 3095 11970 3100
rect 11770 3090 11960 3095
rect 12110 3025 12300 4505
rect 9660 2855 9840 2860
rect 10650 3020 11060 3025
rect 10650 2860 10660 3020
rect 11050 2860 11060 3020
rect 12100 3020 12310 3025
rect 12100 2870 12110 3020
rect 12300 2870 12310 3020
rect 12100 2865 12310 2870
rect 12110 2860 12300 2865
rect 10650 2855 11060 2860
rect 5960 980 5970 1140
rect 6190 1130 6430 1140
rect 7660 1135 7900 1140
rect 6190 990 6270 1130
rect 6410 990 6430 1130
rect 6190 980 6430 990
rect 7650 1130 7900 1135
rect 7650 990 7660 1130
rect 7880 1090 7900 1130
rect 7880 990 7890 1090
rect 7650 985 7890 990
rect 7660 980 7890 985
rect 5960 975 6200 980
rect 2890 -420 3690 -415
rect 1260 -460 1640 -455
rect -610 -540 -470 -535
rect -610 -660 -600 -540
rect -480 -660 -470 -540
rect 1260 -630 1270 -460
rect 1630 -630 1640 -460
rect 1260 -635 1640 -630
rect -610 -665 -470 -660
rect -3030 -1005 -2130 -1000
rect -60 -870 140 -865
rect -6280 -1120 -6180 -1115
rect -6280 -1200 -6270 -1120
rect -6190 -1200 -6180 -1120
rect -6280 -1205 -6180 -1200
rect -6280 -1820 -6220 -1205
rect -60 -1230 -50 -870
rect 130 -1230 140 -870
rect 2890 -990 2900 -420
rect 3680 -990 3690 -420
rect 2890 -995 3690 -990
rect 5350 -430 6050 -425
rect 5350 -1000 5360 -430
rect 6040 -1000 6050 -430
rect 6270 -485 6410 980
rect 6510 895 6650 900
rect 6500 890 6660 895
rect 6500 750 6510 890
rect 6650 750 6660 890
rect 6500 745 6660 750
rect 6260 -490 6420 -485
rect 6260 -630 6270 -490
rect 6410 -630 6420 -490
rect 6260 -635 6420 -630
rect 6270 -640 6410 -635
rect 6510 -725 6650 745
rect 6890 -475 7220 960
rect 6880 -480 7230 -475
rect 6880 -640 6890 -480
rect 7220 -640 7230 -480
rect 7660 -485 7800 980
rect 7890 895 8030 900
rect 7880 890 8040 895
rect 7880 750 7890 890
rect 8030 750 8040 890
rect 7880 745 8040 750
rect 7650 -490 7810 -485
rect 7650 -630 7660 -490
rect 7800 -630 7810 -490
rect 7650 -635 7810 -630
rect 7660 -640 7800 -635
rect 6880 -645 7230 -640
rect 7890 -725 8030 745
rect 8390 -485 8590 2855
rect 10830 1150 11240 1155
rect 9870 1135 10010 1140
rect 9860 1130 10020 1135
rect 9860 990 9870 1130
rect 10010 990 10020 1130
rect 9860 985 10020 990
rect 10830 990 10840 1150
rect 11230 990 11240 1150
rect 11870 1135 12010 1140
rect 10830 985 11240 990
rect 11860 1130 12020 1135
rect 11860 990 11870 1130
rect 12010 990 12020 1130
rect 11860 985 12020 990
rect 9300 -420 9640 -415
rect 8380 -490 8600 -485
rect 8380 -630 8390 -490
rect 8590 -630 8600 -490
rect 8380 -635 8600 -630
rect 6500 -730 6660 -725
rect 6500 -870 6510 -730
rect 6650 -870 6660 -730
rect 6500 -875 6660 -870
rect 7880 -730 8040 -725
rect 7880 -870 7890 -730
rect 8030 -870 8040 -730
rect 7880 -875 8040 -870
rect 6510 -880 6650 -875
rect 7890 -880 8030 -875
rect 5350 -1005 6050 -1000
rect 9300 -1000 9310 -420
rect 9630 -1000 9640 -420
rect 9870 -485 10010 985
rect 10130 895 10270 900
rect 10120 890 10280 895
rect 10120 750 10130 890
rect 10270 750 10280 890
rect 10120 745 10280 750
rect 9860 -490 10020 -485
rect 9860 -630 9870 -490
rect 10010 -630 10020 -490
rect 9860 -635 10020 -630
rect 9870 -640 10010 -635
rect 10130 -725 10270 745
rect 10840 -485 11230 985
rect 11870 -485 12010 985
rect 12160 895 12300 900
rect 12150 890 12310 895
rect 12150 750 12160 890
rect 12300 750 12310 890
rect 12150 745 12310 750
rect 10830 -490 11240 -485
rect 10830 -630 10840 -490
rect 11230 -630 11240 -490
rect 10830 -635 11240 -630
rect 11860 -490 12020 -485
rect 11860 -630 11870 -490
rect 12010 -630 12020 -490
rect 11860 -635 12020 -630
rect 10840 -640 11230 -635
rect 11870 -640 12010 -635
rect 12160 -725 12300 745
rect 10120 -730 10280 -725
rect 10120 -870 10130 -730
rect 10270 -870 10280 -730
rect 10120 -875 10280 -870
rect 12150 -730 12310 -725
rect 12150 -870 12160 -730
rect 12300 -870 12310 -730
rect 12150 -875 12310 -870
rect 10130 -880 10270 -875
rect 12160 -880 12300 -875
rect 9300 -1005 9640 -1000
rect -60 -1235 140 -1230
rect 9020 -1230 9150 -1225
rect 9020 -1350 9030 -1230
rect 9140 -1350 9150 -1230
rect 9020 -1355 9150 -1350
rect 20 -1740 120 -1735
rect -1030 -1800 -950 -1795
rect -1030 -1820 -1020 -1800
rect -6280 -1870 -1020 -1820
rect -960 -1870 -950 -1800
rect 20 -1830 30 -1740
rect 110 -1770 120 -1740
rect 9070 -1770 9130 -1355
rect 110 -1830 9130 -1770
rect 20 -1835 120 -1830
rect -6280 -1875 -950 -1870
rect -6280 -1880 -990 -1875
<< via3 >>
rect -6280 7040 -5770 7560
rect -1200 7060 -570 7530
rect 2990 7070 3620 7540
rect 8470 7080 9100 7550
rect -6850 -1000 -6350 -410
rect -3020 -1000 -2140 -420
rect 1190 2640 1320 3020
rect 1530 3010 1670 3030
rect 1530 2860 1670 3010
rect 1530 2640 1670 2860
rect 1270 -630 1630 -460
rect -50 -1230 130 -870
rect 2900 -990 3680 -420
rect 5360 -1000 6040 -430
rect 9310 -1000 9630 -420
<< metal4 >>
rect -6281 7560 -5769 7561
rect -6281 7040 -6280 7560
rect -5770 7040 -5769 7560
rect 8469 7550 9101 7551
rect 2989 7540 3621 7541
rect -1201 7530 -569 7531
rect -1201 7060 -1200 7530
rect -570 7060 -569 7530
rect 2989 7070 2990 7540
rect 3620 7070 3621 7540
rect 8469 7080 8470 7550
rect 9100 7080 9101 7550
rect 8469 7079 9101 7080
rect 2989 7069 3621 7070
rect -1201 7059 -569 7060
rect -6281 7039 -5769 7040
rect 210 2860 480 3260
rect 1529 3030 1671 3031
rect 1189 3020 1321 3021
rect 630 2640 1190 3020
rect 1320 2640 1321 3020
rect 1189 2639 1321 2640
rect 1529 2640 1530 3030
rect 1670 3010 1671 3030
rect 1670 2640 1671 2660
rect 1529 2639 1671 2640
rect 670 1940 2150 2310
rect -6851 -410 -6349 -409
rect -6851 -1000 -6850 -410
rect -6350 -1000 -6349 -410
rect -6851 -1001 -6349 -1000
rect -3021 -420 -2139 -419
rect -3021 -1000 -3020 -420
rect -2140 -1000 -2139 -420
rect 2899 -420 3681 -419
rect 1269 -460 1631 -459
rect 1269 -630 1270 -460
rect 1630 -630 1631 -460
rect 1269 -631 1631 -630
rect -51 -870 131 -869
rect -3021 -1001 -2139 -1000
rect -1310 -1230 -50 -870
rect 130 -1230 131 -870
rect -51 -1231 131 -1230
rect 1270 -1310 1630 -631
rect 2899 -990 2900 -420
rect 3680 -990 3681 -420
rect 9309 -420 9631 -419
rect 2899 -991 3681 -990
rect 5359 -430 6041 -429
rect 5359 -1000 5360 -430
rect 6040 -1000 6041 -430
rect 5359 -1001 6041 -1000
rect 9309 -1000 9310 -420
rect 9630 -1000 9631 -420
rect 9309 -1001 9631 -1000
rect 700 -1380 2630 -1310
rect 700 -1850 2470 -1380
<< via4 >>
rect -6280 7040 -5770 7560
rect -1200 7060 -570 7530
rect 2990 7070 3620 7540
rect 8470 7080 9100 7550
rect 1530 2660 1670 3010
rect 1670 2660 1860 3010
rect -6850 -1000 -6350 -410
rect -3020 -1000 -2140 -420
rect 2900 -990 3680 -420
rect 5360 -1000 6040 -430
rect 9310 -1000 9630 -420
<< metal5 >>
rect -6304 7570 -5746 7584
rect 4360 7570 5040 7580
rect 8446 7570 9124 7574
rect -9610 7560 12600 7570
rect -9610 7040 -6280 7560
rect -5770 7550 12600 7560
rect -5770 7540 8470 7550
rect -5770 7530 2990 7540
rect -5770 7060 -1200 7530
rect -570 7070 2990 7530
rect 3620 7080 8470 7540
rect 9100 7080 12600 7550
rect 3620 7070 12600 7080
rect -570 7060 12600 7070
rect -5770 7040 12600 7060
rect -9610 6510 -9210 7040
rect -6310 6580 -5740 7040
rect -1224 7036 -546 7040
rect 9910 6550 10340 7040
rect 12040 6480 12600 7040
rect 1500 3010 2310 3040
rect 1500 2660 1530 3010
rect 1860 2660 2310 3010
rect 1500 2630 2310 2660
rect 670 1940 2150 2310
rect -9590 -400 -9160 310
rect -6340 -386 -5590 340
rect -6874 -400 -5590 -386
rect 8790 -396 9340 400
rect -3044 -400 -2116 -396
rect 2876 -400 3704 -396
rect 8790 -400 9654 -396
rect 12200 -400 12750 370
rect -9590 -410 12750 -400
rect -9590 -1000 -6850 -410
rect -6350 -420 12750 -410
rect -6350 -1000 -3020 -420
rect -2140 -990 2900 -420
rect 3680 -430 9310 -420
rect 3680 -990 5360 -430
rect -2140 -1000 5360 -990
rect 6040 -1000 9310 -430
rect 9630 -1000 12750 -420
rect -9590 -1010 12750 -1000
rect -6874 -1024 -6326 -1010
rect -3044 -1024 -2116 -1010
rect -90 -1850 550 -1010
rect 2370 -1014 3704 -1010
rect 2370 -1850 3010 -1014
rect 5336 -1024 6064 -1010
rect 9286 -1024 9654 -1010
use currm_n  currm_n_0
timestamp 1653925904
transform 1 0 820 0 1 590
box -60 -870 658 760
use currm_n  currm_n_1
timestamp 1653925904
transform 1 0 1520 0 1 590
box -60 -870 658 760
use currm_n  currm_n_2
timestamp 1653925904
transform 1 0 2220 0 1 590
box -60 -870 658 760
use currm_n  currm_n_3
timestamp 1653925904
transform 1 0 120 0 1 590
box -60 -870 658 760
use currm_n  currm_n_4
timestamp 1653925904
transform 1 0 2920 0 1 590
box -60 -870 658 760
use currm_n  currm_n_5
timestamp 1653925904
transform 1 0 -580 0 1 590
box -60 -870 658 760
use currm_n  currm_n_6
timestamp 1653925904
transform 1 0 4010 0 1 590
box -60 -870 658 760
use currm_n  currm_n_7
timestamp 1653925904
transform 1 0 4710 0 1 590
box -60 -870 658 760
use currm_n  currm_n_8
timestamp 1653925904
transform 1 0 5410 0 1 590
box -60 -870 658 760
use currm_n  currm_n_9
timestamp 1653925904
transform 1 0 7510 0 1 590
box -60 -870 658 760
use currm_n  currm_n_10
timestamp 1653925904
transform 1 0 6810 0 1 590
box -60 -870 658 760
use currm_n  currm_n_11
timestamp 1653925904
transform 1 0 6110 0 1 590
box -60 -870 658 760
use currm_n  currm_n_12
timestamp 1653925904
transform 1 0 7510 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_13
timestamp 1653925904
transform 1 0 6810 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_14
timestamp 1653925904
transform 1 0 6110 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_15
timestamp 1653925904
transform 1 0 -5170 0 1 590
box -60 -870 658 760
use currm_n  currm_n_16
timestamp 1653925904
transform 1 0 -4470 0 1 590
box -60 -870 658 760
use currm_n  currm_n_17
timestamp 1653925904
transform 1 0 -3770 0 1 590
box -60 -870 658 760
use currm_n  currm_n_18
timestamp 1653925904
transform 1 0 -2370 0 1 590
box -60 -870 658 760
use currm_n  currm_n_19
timestamp 1653925904
transform 1 0 -3070 0 1 590
box -60 -870 658 760
use currm_n  currm_n_20
timestamp 1653925904
transform 1 0 -1670 0 1 590
box -60 -870 658 760
use currm_n  currm_n_21
timestamp 1653925904
transform 1 0 -5170 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_22
timestamp 1653925904
transform 1 0 -3770 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_23
timestamp 1653925904
transform 1 0 -4470 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_24
timestamp 1653925904
transform 1 0 8210 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_25
timestamp 1653925904
transform 1 0 -5870 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_26
timestamp 1653925904
transform 1 0 -6760 0 1 590
box -60 -870 658 760
use currm_n  currm_n_27
timestamp 1653925904
transform 1 0 -8860 0 1 590
box -60 -870 658 760
use currm_n  currm_n_28
timestamp 1653925904
transform 1 0 -8160 0 1 590
box -60 -870 658 760
use currm_n  currm_n_29
timestamp 1653925904
transform 1 0 -7460 0 1 590
box -60 -870 658 760
use currm_n  currm_n_30
timestamp 1653925904
transform 1 0 -9560 0 1 590
box -60 -870 658 760
use currm_n  currm_n_31
timestamp 1653925904
transform 1 0 -9560 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_32
timestamp 1653925904
transform 1 0 11800 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_33
timestamp 1653925904
transform 1 0 -5870 0 1 590
box -60 -870 658 760
use currm_n  currm_n_34
timestamp 1653925904
transform 1 0 -8860 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_35
timestamp 1653925904
transform 1 0 9700 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_36
timestamp 1653925904
transform 1 0 10400 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_37
timestamp 1653925904
transform 1 0 11100 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_38
timestamp 1653925904
transform 1 0 9000 0 1 590
box -60 -870 658 760
use currm_n  currm_n_39
timestamp 1653925904
transform 1 0 11100 0 1 590
box -60 -870 658 760
use currm_n  currm_n_40
timestamp 1653925904
transform 1 0 10400 0 1 590
box -60 -870 658 760
use currm_n  currm_n_41
timestamp 1653925904
transform 1 0 9700 0 1 590
box -60 -870 658 760
use currm_n  currm_n_42
timestamp 1653925904
transform 1 0 11800 0 1 590
box -60 -870 658 760
use currm_n  currm_n_43
timestamp 1653925904
transform 1 0 8210 0 1 590
box -60 -870 658 760
use currm_n  currm_n_44
timestamp 1653925904
transform 1 0 1520 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_45
timestamp 1653925904
transform 1 0 2220 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_46
timestamp 1653925904
transform 1 0 120 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_47
timestamp 1653925904
transform 1 0 820 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_48
timestamp 1653925904
transform 1 0 -8160 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_49
timestamp 1653925904
transform 1 0 -7460 0 1 -1030
box -60 -870 658 760
use currm_p  currm_p_0
timestamp 1653925904
transform 1 0 170 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_1
timestamp 1653925904
transform 1 0 1510 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_2
timestamp 1653925904
transform 1 0 -1170 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_3
timestamp 1653925904
transform 1 0 -2510 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_4
timestamp 1653925904
transform 1 0 -2510 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_5
timestamp 1653925904
transform 1 0 -2510 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_6
timestamp 1653925904
transform 1 0 -3850 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_7
timestamp 1653925904
transform 1 0 -3850 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_8
timestamp 1653925904
transform 1 0 -3850 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_9
timestamp 1653925904
transform 1 0 -5190 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_10
timestamp 1653925904
transform 1 0 -5190 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_11
timestamp 1653925904
transform 1 0 -5190 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_12
timestamp 1653925904
transform 1 0 2850 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_13
timestamp 1653925904
transform 1 0 6870 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_14
timestamp 1653925904
transform 1 0 6870 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_15
timestamp 1653925904
transform 1 0 6870 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_16
timestamp 1653925904
transform 1 0 5530 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_17
timestamp 1653925904
transform 1 0 5530 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_18
timestamp 1653925904
transform 1 0 5530 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_19
timestamp 1653925904
transform 1 0 4190 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_20
timestamp 1653925904
transform 1 0 4190 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_21
timestamp 1653925904
transform 1 0 4190 0 1 3450
box -60 -810 1298 848
use currm_ps  currm_ps_0
timestamp 1653409843
transform 1 0 8200 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_1
timestamp 1653409843
transform 1 0 9290 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_2
timestamp 1653409843
transform 1 0 9290 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_3
timestamp 1653409843
transform 1 0 9290 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_4
timestamp 1653409843
transform 1 0 10380 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_5
timestamp 1653409843
transform 1 0 10380 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_6
timestamp 1653409843
transform 1 0 10380 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_7
timestamp 1653409843
transform 1 0 11470 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_8
timestamp 1653409843
transform 1 0 11470 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_9
timestamp 1653409843
transform 1 0 11470 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_10
timestamp 1653409843
transform 1 0 8200 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_11
timestamp 1653409843
transform 1 0 -7380 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_12
timestamp 1653409843
transform 1 0 -9560 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_13
timestamp 1653409843
transform 1 0 -8470 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_14
timestamp 1653409843
transform 1 0 -7380 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_15
timestamp 1653409843
transform 1 0 -7380 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_16
timestamp 1653409843
transform 1 0 -9560 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_17
timestamp 1653409843
transform 1 0 -8470 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_18
timestamp 1653409843
transform 1 0 -6290 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_19
timestamp 1653409843
transform 1 0 -6290 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_20
timestamp 1653409843
transform 1 0 -9560 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_21
timestamp 1653409843
transform 1 0 -8470 0 1 2690
box -50 -50 1052 1608
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_2
timestamp 1653925904
transform 0 1 -2159 -1 0 3473
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_3
timestamp 1653925904
transform 0 1 5041 -1 0 3483
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_MJMGTW  sky130_fd_pr__cap_mim_m3_2_MJMGTW_0
timestamp 1653911185
transform 0 1 10711 -1 0 3483
box -3351 -2101 3373 2101
use sky130_fd_pr__cap_mim_m3_2_MJMGTW  sky130_fd_pr__cap_mim_m3_2_MJMGTW_1
timestamp 1653911185
transform 0 1 -7689 -1 0 3443
box -3351 -2101 3373 2101
use sky130_fd_pr__cap_mim_m3_2_N3PKNJ  sky130_fd_pr__cap_mim_m3_2_N3PKNJ_0
timestamp 1653911185
transform 1 0 -2149 0 1 -2449
box -3351 -1101 3373 1101
use sky130_fd_pr__cap_mim_m3_2_N3PKNJ  sky130_fd_pr__cap_mim_m3_2_N3PKNJ_1
timestamp 1653911185
transform -1 0 5083 0 -1 -2449
box -3351 -1101 3373 1101
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_0
timestamp 1653899151
transform 1 0 -669 0 1 -1560
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_E6B2KN  sky130_fd_pr__nfet_01v8_E6B2KN_0
timestamp 1653925904
transform 1 0 1155 0 1 1760
box -325 -410 325 410
use sky130_fd_pr__nfet_01v8_E6B2KN  sky130_fd_pr__nfet_01v8_E6B2KN_1
timestamp 1653925904
transform 1 0 1795 0 1 1760
box -325 -410 325 410
use sky130_fd_pr__nfet_01v8_LH2JGW  sky130_fd_pr__nfet_01v8_LH2JGW_0
timestamp 1653925904
transform 1 0 -207 0 1 -1460
box -263 -410 263 410
use sky130_fd_pr__nfet_01v8_LH2JGW  sky130_fd_pr__nfet_01v8_LH2JGW_1
timestamp 1653925904
transform 1 0 -6177 0 1 -680
box -263 -410 263 410
use sky130_fd_pr__nfet_01v8_LH2JGW  sky130_fd_pr__nfet_01v8_LH2JGW_2
timestamp 1653925904
transform 1 0 9123 0 1 -690
box -263 -410 263 410
use sky130_fd_pr__pfet_01v8_U47ZGH  sky130_fd_pr__pfet_01v8_U47ZGH_0
timestamp 1653925904
transform 1 0 -5981 0 1 6339
box -359 -419 359 419
use sky130_fd_pr__pfet_01v8_U47ZGH  sky130_fd_pr__pfet_01v8_U47ZGH_1
timestamp 1653925904
transform 1 0 8509 0 1 6339
box -359 -419 359 419
use sky130_fd_pr__pfet_01v8_UAQRRG  sky130_fd_pr__pfet_01v8_UAQRRG_0
timestamp 1653899151
transform 1 0 -689 0 1 -911
box -211 -319 211 319
<< labels >>
rlabel metal2 1440 -640 1490 -540 1 I_Bias
rlabel metal1 -490 -1740 -440 -1690 1 Disable_FB
rlabel metal1 1310 1990 1390 2060 1 InP
rlabel metal1 1540 1990 1620 2060 1 InN
rlabel metal5 -6580 7180 -6380 7500 1 VP
rlabel metal2 11820 1690 12190 2060 1 OutN
rlabel metal3 -7670 1780 -7300 2150 1 OutP
rlabel metal5 4080 -920 4600 -540 1 VN
rlabel metal1 -820 -380 -790 -350 1 Disable_FB_B
rlabel metal3 7710 1770 7880 1960 1 VM34D
rlabel metal1 9000 1390 9030 1420 1 VM31D
rlabel metal1 -6320 1590 -6290 1630 1 VM30D
rlabel space -4970 1880 -4770 2080 1 VM9D
rlabel metal2 990 2420 1170 2500 1 VM16D
rlabel metal2 1770 2410 1950 2490 1 VM14D
<< end >>
