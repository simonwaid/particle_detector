magic
tech sky130A
magscale 1 2
timestamp 1646301356
<< pwell >>
rect -5618 -998 5618 998
<< psubdiff >>
rect -5582 928 -5486 962
rect 5486 928 5582 962
rect -5582 866 -5548 928
rect 5548 866 5582 928
rect -5582 -928 -5548 -866
rect 5548 -928 5582 -866
rect -5582 -962 -5486 -928
rect 5486 -962 5582 -928
<< psubdiffcont >>
rect -5486 928 5486 962
rect -5582 -866 -5548 866
rect 5548 -866 5582 866
rect -5486 -962 5486 -928
<< xpolycontact >>
rect -5452 400 -4306 832
rect -5452 -832 -4306 -400
rect -4058 400 -2912 832
rect -4058 -832 -2912 -400
rect -2664 400 -1518 832
rect -2664 -832 -1518 -400
rect -1270 400 -124 832
rect -1270 -832 -124 -400
rect 124 400 1270 832
rect 124 -832 1270 -400
rect 1518 400 2664 832
rect 1518 -832 2664 -400
rect 2912 400 4058 832
rect 2912 -832 4058 -400
rect 4306 400 5452 832
rect 4306 -832 5452 -400
<< ppolyres >>
rect -5452 -400 -4306 400
rect -4058 -400 -2912 400
rect -2664 -400 -1518 400
rect -1270 -400 -124 400
rect 124 -400 1270 400
rect 1518 -400 2664 400
rect 2912 -400 4058 400
rect 4306 -400 5452 400
<< locali >>
rect -5582 928 -5486 962
rect 5486 928 5582 962
rect -5582 866 -5548 928
rect 5548 866 5582 928
rect -5582 -928 -5548 -866
rect 5548 -928 5582 -866
rect -5582 -962 -5486 -928
rect 5486 -962 5582 -928
<< viali >>
rect -5436 417 -4322 814
rect -4042 417 -2928 814
rect -2648 417 -1534 814
rect -1254 417 -140 814
rect 140 417 1254 814
rect 1534 417 2648 814
rect 2928 417 4042 814
rect 4322 417 5436 814
rect -5436 -814 -4322 -417
rect -4042 -814 -2928 -417
rect -2648 -814 -1534 -417
rect -1254 -814 -140 -417
rect 140 -814 1254 -417
rect 1534 -814 2648 -417
rect 2928 -814 4042 -417
rect 4322 -814 5436 -417
<< metal1 >>
rect -5448 814 -4310 820
rect -5448 417 -5436 814
rect -4322 417 -4310 814
rect -5448 411 -4310 417
rect -4054 814 -2916 820
rect -4054 417 -4042 814
rect -2928 417 -2916 814
rect -4054 411 -2916 417
rect -2660 814 -1522 820
rect -2660 417 -2648 814
rect -1534 417 -1522 814
rect -2660 411 -1522 417
rect -1266 814 -128 820
rect -1266 417 -1254 814
rect -140 417 -128 814
rect -1266 411 -128 417
rect 128 814 1266 820
rect 128 417 140 814
rect 1254 417 1266 814
rect 128 411 1266 417
rect 1522 814 2660 820
rect 1522 417 1534 814
rect 2648 417 2660 814
rect 1522 411 2660 417
rect 2916 814 4054 820
rect 2916 417 2928 814
rect 4042 417 4054 814
rect 2916 411 4054 417
rect 4310 814 5448 820
rect 4310 417 4322 814
rect 5436 417 5448 814
rect 4310 411 5448 417
rect -5448 -417 -4310 -411
rect -5448 -814 -5436 -417
rect -4322 -814 -4310 -417
rect -5448 -820 -4310 -814
rect -4054 -417 -2916 -411
rect -4054 -814 -4042 -417
rect -2928 -814 -2916 -417
rect -4054 -820 -2916 -814
rect -2660 -417 -1522 -411
rect -2660 -814 -2648 -417
rect -1534 -814 -1522 -417
rect -2660 -820 -1522 -814
rect -1266 -417 -128 -411
rect -1266 -814 -1254 -417
rect -140 -814 -128 -417
rect -1266 -820 -128 -814
rect 128 -417 1266 -411
rect 128 -814 140 -417
rect 1254 -814 1266 -417
rect 128 -820 1266 -814
rect 1522 -417 2660 -411
rect 1522 -814 1534 -417
rect 2648 -814 2660 -417
rect 1522 -820 2660 -814
rect 2916 -417 4054 -411
rect 2916 -814 2928 -417
rect 4042 -814 4054 -417
rect 2916 -820 4054 -814
rect 4310 -417 5448 -411
rect 4310 -814 4322 -417
rect 5436 -814 5448 -417
rect 4310 -820 5448 -814
<< res5p73 >>
rect -5454 -402 -4304 402
rect -4060 -402 -2910 402
rect -2666 -402 -1516 402
rect -1272 -402 -122 402
rect 122 -402 1272 402
rect 1516 -402 2666 402
rect 2910 -402 4060 402
rect 4304 -402 5454 402
<< properties >>
string FIXED_BBOX -5565 -945 5565 945
string gencell sky130_fd_pr__res_high_po_5p73
string library sky130
string parameters w 5.730 l 4 m 1 nx 8 wmin 5.730 lmin 0.50 rho 319.8 val 291.246 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 5.730 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
