magic
tech sky130A
magscale 1 2
timestamp 1645462850
<< pwell >>
rect -307 -1598 307 1598
<< psubdiff >>
rect -271 1528 -175 1562
rect 175 1528 271 1562
rect -271 1466 -237 1528
rect 237 1466 271 1528
rect -271 -1528 -237 -1466
rect 237 -1528 271 -1466
rect -271 -1562 -175 -1528
rect 175 -1562 271 -1528
<< psubdiffcont >>
rect -175 1528 175 1562
rect -271 -1466 -237 1466
rect 237 -1466 271 1466
rect -175 -1562 175 -1528
<< xpolycontact >>
rect -141 1000 141 1432
rect -141 -1432 141 -1000
<< xpolyres >>
rect -141 -1000 141 1000
<< locali >>
rect -271 1528 -175 1562
rect 175 1528 271 1562
rect -271 1466 -237 1528
rect 237 1466 271 1528
rect -271 -1528 -237 -1466
rect 237 -1528 271 -1466
rect -271 -1562 -175 -1528
rect 175 -1562 271 -1528
<< viali >>
rect -125 1017 125 1414
rect -125 -1414 125 -1017
<< metal1 >>
rect -131 1414 131 1426
rect -131 1017 -125 1414
rect 125 1017 131 1414
rect -131 1005 131 1017
rect -131 -1017 131 -1005
rect -131 -1414 -125 -1017
rect 125 -1414 131 -1017
rect -131 -1426 131 -1414
<< res1p41 >>
rect -143 -1002 143 1002
<< properties >>
string FIXED_BBOX -254 -1545 254 1545
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 10 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 14.451k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
