magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< dnwell >>
rect 70 8020 3300 9920
<< nwell >>
rect -10 9714 3380 10000
rect -10 8226 276 9714
rect 3094 8226 3380 9714
rect -10 7940 3380 8226
<< pwell >>
rect 276 8226 3094 9714
<< nsubdiff >>
rect 27 9943 3343 9963
rect 27 9909 107 9943
rect 3263 9909 3343 9943
rect 27 9889 3343 9909
rect 27 9883 101 9889
rect 27 8057 47 9883
rect 81 8057 101 9883
rect 27 8051 101 8057
rect 3269 9883 3343 9889
rect 3269 8057 3289 9883
rect 3323 8057 3343 9883
rect 3269 8051 3343 8057
rect 27 8031 3343 8051
rect 27 7997 107 8031
rect 3263 7997 3343 8031
rect 27 7977 3343 7997
<< nsubdiffcont >>
rect 107 9909 3263 9943
rect 47 8057 81 9883
rect 3289 8057 3323 9883
rect 107 7997 3263 8031
<< locali >>
rect 1640 11620 1730 12370
rect 1630 10090 1750 11620
rect -520 7690 -310 10070
rect 1640 10050 1740 10090
rect 20 9950 3340 9960
rect 20 9943 1600 9950
rect 1790 9943 3340 9950
rect 20 9909 107 9943
rect 3263 9909 3340 9943
rect 20 9890 1600 9909
rect 20 9883 100 9890
rect 20 8057 47 9883
rect 81 8057 100 9883
rect 1790 9890 3340 9909
rect 3270 9883 3340 9890
rect 1620 9240 1750 9650
rect 1620 8290 1750 8700
rect 20 8050 100 8057
rect 3270 8057 3289 9883
rect 3323 8057 3340 9883
rect 3270 8050 3340 8057
rect 20 8031 3340 8050
rect 20 7997 107 8031
rect 3263 7997 3340 8031
rect 20 7980 3340 7997
rect 3530 7690 3740 10070
rect -520 7520 10 7690
rect 1840 7520 3740 7690
rect 2800 120 3290 7520
rect 930 -190 3290 120
rect 930 -280 980 -190
rect 1940 -280 3290 -190
<< viali >>
rect 1600 9943 1790 9950
rect 1600 9909 1790 9943
rect 1600 9840 1790 9909
rect 1620 8700 1750 9240
rect 980 -280 1940 -190
<< metal1 >>
rect -1510 11800 4870 12250
rect -1500 10180 -1490 10620
rect 1530 10180 1540 10620
rect 1600 9956 1790 11800
rect 1830 10170 1840 10620
rect 4870 10170 4880 10620
rect 1588 9950 1802 9956
rect 1588 9840 1600 9950
rect 1790 9840 1802 9950
rect 1588 9834 1802 9840
rect 310 9510 1510 9590
rect 1860 9510 3060 9590
rect 310 9050 390 9510
rect 1614 9240 1756 9252
rect 310 9040 1510 9050
rect 260 8900 270 9040
rect 380 8900 1510 9040
rect 310 8890 1510 8900
rect 310 8430 390 8890
rect 1610 8700 1620 9240
rect 1750 8700 1760 9240
rect 2980 9050 3060 9510
rect 1860 9040 3060 9050
rect 1860 8900 2990 9040
rect 3100 8900 3110 9040
rect 1860 8890 3060 8900
rect 1614 8688 1756 8700
rect 2980 8430 3060 8890
rect 310 8350 1510 8430
rect 1860 8350 3060 8430
rect 968 -190 1952 -184
rect 968 -280 980 -190
rect 1940 -280 1952 -190
rect 968 -286 1952 -280
<< via1 >>
rect -1490 10180 1530 10620
rect 1840 10170 4870 10620
rect 270 8900 380 9040
rect 1620 8700 1750 9240
rect 2990 8900 3100 9040
rect 980 -280 1940 -190
<< metal2 >>
rect -1490 10620 1530 10630
rect -1490 10170 450 10180
rect 990 10170 1530 10180
rect 1840 10620 4870 10630
rect 450 10160 990 10170
rect 1840 10160 4870 10170
rect -1610 9620 3060 9750
rect 260 9040 390 9620
rect 440 9470 1450 9480
rect 440 9330 450 9470
rect 980 9330 1450 9470
rect 440 9320 1450 9330
rect 1910 9470 2920 9480
rect 1910 9330 2380 9470
rect 2910 9330 2920 9470
rect 1910 9320 2920 9330
rect 1620 9240 1750 9250
rect 530 9230 1620 9240
rect 1750 9230 2830 9240
rect 530 9090 1090 9230
rect 2280 9090 2830 9230
rect 530 9080 1620 9090
rect 260 8900 270 9040
rect 380 8900 390 9040
rect 260 8890 390 8900
rect 530 8850 1620 8860
rect 1750 9080 2830 9090
rect 2980 9040 3110 9050
rect 2980 8900 2990 9040
rect 3100 8900 3110 9040
rect 1750 8850 2830 8860
rect 530 8710 1090 8850
rect 2280 8710 2830 8850
rect 530 8700 1620 8710
rect 1750 8700 2830 8710
rect 1620 8690 1750 8700
rect 440 8610 1450 8620
rect 440 8470 450 8610
rect 980 8470 1450 8610
rect 440 8460 1450 8470
rect 1910 8610 2920 8620
rect 1910 8470 2380 8610
rect 2910 8470 2920 8610
rect 1910 8460 2920 8470
rect 2980 8190 3110 8900
rect -1610 8060 3110 8190
rect 980 120 1940 130
rect 980 -290 1940 -280
<< via2 >>
rect 450 10180 990 10620
rect 450 10170 990 10180
rect 2370 10170 2910 10620
rect 450 9330 980 9470
rect 2380 9330 2910 9470
rect 1090 9090 1620 9230
rect 1620 9090 1750 9230
rect 1750 9090 2280 9230
rect 1090 8710 1620 8850
rect 1620 8710 1750 8850
rect 1750 8710 2280 8850
rect 450 8470 980 8610
rect 2380 8470 2910 8610
rect 980 -190 1940 120
rect 980 -280 1940 -190
<< metal3 >>
rect 440 10620 1000 10625
rect 440 10170 450 10620
rect 990 10170 1000 10620
rect 440 10165 1000 10170
rect 2360 10620 2920 10625
rect 2360 10170 2370 10620
rect 2910 10170 2920 10620
rect 2360 10165 2920 10170
rect 440 9980 990 10165
rect 440 9600 450 9980
rect 980 9600 990 9980
rect 440 9470 990 9600
rect 440 9330 450 9470
rect 980 9330 990 9470
rect 440 8610 990 9330
rect 2370 9470 2920 10165
rect 2370 9330 2380 9470
rect 2910 9330 2920 9470
rect 440 8470 450 8610
rect 980 8470 990 8610
rect 440 8460 990 8470
rect 1080 9230 2290 9240
rect 1080 9090 1090 9230
rect 2280 9090 2290 9230
rect 1080 8850 2290 9090
rect 1080 8710 1090 8850
rect 2280 8710 2290 8850
rect 1080 8160 2290 8710
rect 2370 8610 2920 9330
rect 2370 8470 2380 8610
rect 2910 8470 2920 8610
rect 2370 8460 2920 8470
rect 980 8080 2290 8160
rect 980 7910 1720 8080
rect 990 140 1880 650
rect -20 120 2850 140
rect -20 -280 980 120
rect 1940 -280 2850 120
rect -20 -880 2850 -280
<< via3 >>
rect 2380 10210 2910 10590
rect 450 9600 980 9980
<< metal4 >>
rect 440 10590 5040 10600
rect 440 10210 2380 10590
rect 2910 10210 5040 10590
rect 440 10200 5040 10210
rect 440 9980 5040 9990
rect 440 9600 450 9980
rect 980 9600 5040 9980
rect 440 9590 5040 9600
use outd_cmirror_64t  outd_cmirror_64t_0
timestamp 1654768133
transform 1 0 -10 0 1 76
box 0 -76 2862 7840
use outd_diffamp  outd_diffamp_0
timestamp 1654768133
transform 1 0 300 0 1 320
box 0 7930 2768 9368
use sky130_fd_pr__res_high_po_2p85_8GE2XM  sky130_fd_pr__res_high_po_2p85_8GE2XM_0
timestamp 1654768133
transform 1 0 18 0 1 11208
box -1678 -1198 1678 1198
use sky130_fd_pr__res_high_po_2p85_8GE2XM  sky130_fd_pr__res_high_po_2p85_8GE2XM_1
timestamp 1654768133
transform 1 0 3358 0 1 11208
box -1678 -1198 1678 1198
<< labels >>
rlabel metal3 420 -570 630 -300 1 VN
rlabel metal3 1630 8200 1730 8310 1 isource_out
<< end >>
