* SPICE3 file created from outd.ext - technology: sky130A

X0 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2 VN I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 VN I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X4 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5 VP V_da2_N VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6 VP V_da2_P VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7 V_da2_N VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8 V_da2_P VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9 VP V_da2_P VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10 VP V_da2_N VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11 V_da2_N VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12 VP V_da2_P VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13 V_da2_P VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14 VP V_da2_N VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X15 V_da2_N VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X16 V_da2_P VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X17 VP V_da2_P VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X18 VP V_da2_N VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X19 V_da2_N VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X20 V_da2_P VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X21 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X39 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X40 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X41 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X42 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X43 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X45 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X48 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X51 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X53 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X56 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X57 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X58 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X59 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X61 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X64 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X65 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X66 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X67 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X69 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X70 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X72 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X75 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X76 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X77 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X80 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X83 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X85 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X90 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X92 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X93 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X94 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X98 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X99 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X100 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X101 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X102 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X104 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X105 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X106 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X107 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X108 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X109 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X110 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X111 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X112 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X113 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X114 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X115 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X116 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X117 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X118 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X119 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X120 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X121 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X122 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X123 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X124 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X125 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X126 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X127 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X128 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X129 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X130 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X131 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X132 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X133 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X134 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X135 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X136 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X137 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X138 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X139 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X140 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X141 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X142 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X143 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X145 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X146 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X147 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X148 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X149 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X150 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X151 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X152 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X153 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X154 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X155 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X156 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X157 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X158 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X159 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X160 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X161 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X162 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X163 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X164 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X165 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X166 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X167 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X168 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X169 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X170 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X171 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X172 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X173 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X174 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X175 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X176 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X177 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X178 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X179 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X180 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X181 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X182 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X183 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X184 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X185 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X186 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X187 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X188 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X189 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X190 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X191 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X192 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X193 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X194 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X195 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X196 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X197 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X198 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X199 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X200 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X201 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X202 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X203 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X204 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X205 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X206 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X207 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X208 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X209 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X210 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X211 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X212 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X213 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X214 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X215 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X216 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X217 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X218 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X219 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X220 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X221 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X222 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X223 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X224 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X225 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X226 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X227 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X228 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X229 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X230 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X231 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X232 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X233 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X234 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X235 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X236 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X237 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X238 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X239 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X240 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X241 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X242 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X243 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X244 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X245 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X246 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X247 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X248 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X249 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X250 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X251 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X252 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X253 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X254 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X255 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X256 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X257 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X258 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X259 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X261 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X262 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X263 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X264 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X265 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X266 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X267 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X268 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X269 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X273 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X274 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X275 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X276 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X277 outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X279 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X280 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X281 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X283 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X284 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X285 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X286 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X287 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X288 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X289 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X290 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X291 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X292 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X293 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X294 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X295 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X296 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X297 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X298 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X299 outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X300 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X301 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X302 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X303 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X304 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X305 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X306 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X307 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X308 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X309 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X310 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X311 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X312 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X313 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X314 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X315 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X316 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X317 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X318 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X319 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X320 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X321 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X322 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X323 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X324 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X325 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X326 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X327 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X328 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X329 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X330 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X331 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X332 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X333 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X334 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X335 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X336 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X337 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X338 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X339 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X340 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X341 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X342 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X343 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X344 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X345 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X346 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X347 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X348 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X349 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X350 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X351 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X352 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X353 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X354 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X355 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X356 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X357 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X358 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X359 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X360 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X361 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X362 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X363 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X364 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X365 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X366 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X367 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X368 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X369 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X370 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X371 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X372 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X373 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X374 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X375 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X376 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X377 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X378 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X379 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X380 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X381 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X382 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X383 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X384 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X385 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X386 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X387 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X388 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X389 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X390 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X391 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X392 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X393 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X394 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X395 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X396 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X397 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X398 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X399 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X400 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X401 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X402 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X403 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X404 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X405 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X406 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X407 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X408 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X409 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X410 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X411 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X412 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X413 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X414 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X415 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X416 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X417 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X418 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X419 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X420 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X421 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X422 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X423 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X424 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X425 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X426 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X427 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X428 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X429 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X430 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X431 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X432 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X433 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X434 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X435 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X436 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X437 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X438 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X439 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X440 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X441 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X442 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X443 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X444 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X445 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X446 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X447 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X448 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X449 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X450 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X451 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X452 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X453 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X454 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X455 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X456 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X457 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X458 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X459 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X460 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X461 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X462 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X463 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X464 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X465 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X466 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X467 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X468 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X469 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X470 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X471 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X472 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X473 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X474 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X475 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X476 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X477 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X478 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X479 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X480 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X481 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X482 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X483 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X484 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X485 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X486 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X487 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X488 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X489 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X490 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X491 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X492 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X493 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X494 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X495 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X496 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X497 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X498 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X499 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X500 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X501 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X502 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X503 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X504 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X505 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X506 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X507 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X508 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X509 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X510 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X511 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X512 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X513 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X514 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X515 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X516 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X517 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X519 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X520 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X521 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X522 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X523 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X524 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X525 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X526 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X527 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X528 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X529 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X530 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X531 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X532 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X533 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X534 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X535 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X536 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X537 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X538 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X540 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X541 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X542 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X543 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X544 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X545 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X546 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X547 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X548 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X549 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X550 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X551 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X552 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X553 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X554 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X555 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X556 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X557 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X558 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X559 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X560 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X561 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X562 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X563 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X564 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X565 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X566 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X567 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X568 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X569 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X570 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X571 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X572 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X573 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X574 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X575 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X576 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X577 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X578 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X579 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X580 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X581 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X582 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X583 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X584 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X585 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X586 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X587 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X588 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X589 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X590 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X591 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X592 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X593 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X594 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X595 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X596 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X597 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X598 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X599 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X600 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X601 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X602 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X603 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X604 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X605 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X606 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X607 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X608 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X609 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X610 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X611 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X612 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X613 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X614 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X615 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X616 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X617 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X618 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X619 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X620 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X621 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X622 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X623 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X624 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X625 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X626 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X627 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X628 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X629 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X630 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X631 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X632 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X633 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X634 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X635 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X636 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X637 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X638 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X639 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X640 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X641 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X642 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X643 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X644 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X645 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X646 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X647 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X648 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X649 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X650 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X651 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X652 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X653 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X654 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X655 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X656 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X657 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X658 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X659 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X660 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X661 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X662 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X663 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X664 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X665 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X666 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X667 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X668 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X669 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X670 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X671 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X672 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X673 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X674 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X675 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X676 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X677 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X678 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X679 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X680 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X681 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X682 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X683 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X684 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X685 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X686 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X687 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X688 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X689 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X690 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X691 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X692 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X693 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X694 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X695 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X696 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X697 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X698 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X699 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X700 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X701 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X702 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X703 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X704 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X705 outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X706 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X707 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X708 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X709 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X710 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X711 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X712 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X713 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X714 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X715 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X716 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X717 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X718 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X719 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X720 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X721 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X722 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X723 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X724 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X725 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X726 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X727 outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da1_P V_da2_P outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X728 V_da2_P V_da1_P outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X729 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X730 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X731 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X732 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X733 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X734 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X735 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X736 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X737 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X738 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X739 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X740 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X741 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X742 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X743 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X744 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X745 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X746 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X747 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X748 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X749 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X750 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X751 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X752 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X753 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X754 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X755 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X756 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X757 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X758 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X759 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X760 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X761 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X762 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X763 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X764 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X765 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X766 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X767 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X768 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X769 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X770 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X771 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X772 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X773 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X774 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X775 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X776 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X777 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X778 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X779 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X780 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X781 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X782 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X783 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X784 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X785 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X786 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X787 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X788 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X789 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X790 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X791 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X792 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X793 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X794 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X795 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X796 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X797 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X798 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X799 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X800 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X801 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X802 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X803 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X804 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X805 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X806 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X807 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X808 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X809 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X810 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X811 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X812 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X813 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X814 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X815 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X816 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X817 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X818 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X819 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X820 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X821 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X822 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X823 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X824 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X825 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X826 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X827 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X828 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X829 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X830 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X831 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X832 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X833 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X834 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X835 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X836 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X837 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X838 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X839 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X840 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X841 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X842 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X843 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X844 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X845 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X846 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X847 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X848 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X849 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X850 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X851 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X852 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X853 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X854 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X855 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X856 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X857 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X858 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X859 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X860 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X861 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X862 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X863 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X864 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X865 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X866 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X867 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X868 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X869 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X870 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X871 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X872 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X873 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X874 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X875 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X876 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X877 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X878 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X879 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X880 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X881 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X882 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X883 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X884 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X885 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X886 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X887 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X888 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X889 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X890 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X891 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X892 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X893 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X894 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X895 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X896 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X897 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X898 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X899 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X900 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X901 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X902 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X903 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X904 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X905 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X906 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X907 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X908 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X909 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X910 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X911 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X912 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X913 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X914 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X915 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X916 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X917 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X918 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X919 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X920 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X921 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X922 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X923 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X924 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X925 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X926 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X927 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X928 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X929 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X930 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X931 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X932 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X933 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X934 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X935 VN V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X936 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X937 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X938 VN V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X939 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X940 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X941 outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da1_N V_da2_N outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X942 V_da2_N V_da1_N outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X943 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X944 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X945 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X946 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X947 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X948 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X949 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X950 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X951 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X952 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X953 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X954 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X955 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X956 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X957 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X958 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X959 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X960 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X961 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X962 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X963 VN V_da1_P V_da2_P outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X964 V_da2_P V_da1_P VN outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X965 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X966 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X967 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X968 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X969 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X970 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X971 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X972 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X973 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X974 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X975 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X976 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X977 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X978 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X979 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X980 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X981 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X982 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X983 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X984 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X985 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X986 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X987 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X988 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X989 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X990 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X991 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X992 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X993 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X994 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X995 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X996 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X997 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X998 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X999 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1000 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1001 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1002 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1003 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1004 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1005 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1006 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1007 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1008 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1009 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1010 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1011 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1012 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1013 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1014 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1015 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1016 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1017 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1018 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1019 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1020 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1021 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1022 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1023 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1024 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1025 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1026 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1027 VM1_D I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1028 outd_stage2_0/m2_7240_7300# I_Bias VM1_D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1029 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1030 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1031 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1032 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1033 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1034 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1035 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1036 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1037 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1038 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1039 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1040 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1041 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1042 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1043 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1044 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1045 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1046 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1047 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1048 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1049 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1050 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1051 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1052 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1053 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1054 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1055 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1056 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1057 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1058 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1059 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1060 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1061 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1062 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1063 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1064 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1065 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1066 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1067 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1068 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1069 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1070 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1071 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1072 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1073 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1074 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1075 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1076 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1077 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1078 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1079 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1080 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1081 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1082 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1083 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1084 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1085 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1086 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1087 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1088 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1089 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1090 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1091 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1092 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1093 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1094 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1095 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1096 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1097 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1098 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1099 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1100 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1101 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1102 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1103 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1104 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1105 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1106 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1107 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1108 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1109 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1110 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1111 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1112 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1113 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1114 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1115 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1116 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1117 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1118 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1119 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1120 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1121 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1122 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1123 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1124 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1125 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1126 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1127 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1128 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1129 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1130 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1131 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1132 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1133 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1134 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1135 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1136 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1137 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1138 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1139 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1140 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1141 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1142 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1143 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1144 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1145 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1146 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1147 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1148 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1149 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1150 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1151 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1152 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1153 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1154 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1155 VN I_Bias outd_stage2_0/m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1156 outd_stage2_0/m2_7240_7300# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1157 InputRef VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1158 VN I_Bias m1_n19890_7120# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1159 m1_n19890_7120# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1160 VN I_Bias m1_n19890_7120# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1161 m1_n19890_7120# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1162 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1163 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1164 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1165 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1166 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1167 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1168 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1169 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1170 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1171 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1172 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1173 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1174 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1175 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1176 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1177 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1178 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1179 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1180 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1181 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1182 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1183 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1184 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1185 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1186 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1187 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1188 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1189 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1190 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1191 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1192 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1193 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1194 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1195 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1196 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1197 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1198 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1199 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1200 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1201 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1202 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1203 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1204 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1205 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1206 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1207 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1208 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1209 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1210 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1211 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1212 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1213 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1214 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1215 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1216 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1217 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1218 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1219 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1220 outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1221 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1222 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1223 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1224 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1225 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1226 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1227 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1228 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1229 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1230 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1231 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1232 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1233 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1234 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1235 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1236 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1237 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1238 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1239 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1240 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1241 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1242 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1243 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1244 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1245 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1246 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1247 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1248 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1249 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1250 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1251 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1252 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1253 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1254 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1255 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1256 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1257 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1258 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1259 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1260 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1261 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1262 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1263 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1264 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1265 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1266 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1267 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1268 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1269 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1270 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1271 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1272 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1273 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1274 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1275 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1276 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1277 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1278 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1279 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1280 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1281 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1282 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1283 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1284 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1285 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1286 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1287 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1288 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1289 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1290 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1291 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1292 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1293 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1294 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1295 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1296 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1297 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1298 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1299 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1300 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1301 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1302 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1303 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1304 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1305 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1306 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1307 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1308 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1309 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1310 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1311 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1312 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1313 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1314 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1315 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1316 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1317 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1318 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1319 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1320 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1321 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1322 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1323 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1324 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1325 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1326 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1327 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1328 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1329 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1330 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1331 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1332 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1333 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1334 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1335 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1336 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1337 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1338 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1339 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1340 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1341 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1342 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1343 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1344 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1345 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1346 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1347 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1348 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1349 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1350 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1351 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1352 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1353 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1354 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1355 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1356 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1357 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1358 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1359 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1360 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1361 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1362 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1363 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1364 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1365 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1366 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1367 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1368 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1369 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1370 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1371 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1372 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1373 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1374 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1375 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1376 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1377 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1378 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1379 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1380 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1381 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1382 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1383 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1384 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1385 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1386 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1387 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1388 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1389 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1390 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1391 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1392 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1393 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1394 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1395 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1396 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1397 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1398 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1399 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1400 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1401 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1402 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1403 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1404 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1405 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1406 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1407 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1408 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1409 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1410 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1411 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1412 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1413 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1414 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1415 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1416 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1417 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1418 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1419 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1420 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1421 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1422 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1423 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1424 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1425 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1426 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1427 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1428 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1429 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1430 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1431 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1432 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1433 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1434 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1435 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1436 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1437 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1438 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1439 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1440 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1441 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1442 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1443 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1444 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1445 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1446 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1447 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1448 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1449 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1450 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1451 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1452 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1453 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1454 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1455 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1456 outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1457 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1458 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1459 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1460 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1461 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1462 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1463 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1464 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1465 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1466 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1467 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1468 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1469 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1470 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1471 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1472 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1473 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1474 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1475 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1476 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1477 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1478 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1479 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1480 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1481 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1482 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1483 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1484 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1485 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1486 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1487 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1488 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1489 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1490 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1491 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1492 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1493 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1494 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1495 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1496 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1497 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1498 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1499 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1500 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1501 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1502 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1503 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1504 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1505 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1506 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1507 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1508 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1509 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1510 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1511 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1512 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1513 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1514 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1515 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1516 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1517 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1518 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1519 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1520 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1521 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1522 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1523 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1524 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1525 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1526 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1527 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1528 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1529 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1530 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1531 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1532 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1533 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1534 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1535 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1536 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1537 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1538 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1539 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1540 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1541 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1542 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1543 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1544 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1545 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1546 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1547 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1548 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1549 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1550 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1551 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1552 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1553 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1554 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1555 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1556 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1557 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1558 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1559 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1560 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1561 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1562 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1563 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1564 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1565 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1566 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1567 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1568 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1569 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1570 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1571 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1572 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1573 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1574 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1575 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1576 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1577 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1578 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1579 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1580 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1581 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1582 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1583 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1584 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1585 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1586 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1587 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1588 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1589 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1590 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1591 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1592 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1593 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1594 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1595 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1596 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1597 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1598 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1599 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1600 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1601 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1602 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1603 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1604 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1605 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1606 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1607 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1608 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1609 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1610 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1611 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1612 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1613 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1614 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1615 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1616 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1617 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1618 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1619 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1620 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1621 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1622 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1623 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1624 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1625 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1626 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1627 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1628 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1629 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1630 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1631 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1632 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1633 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1634 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1635 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1636 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1637 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1638 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1639 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1640 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1641 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1642 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1643 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1644 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1645 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1646 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1647 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1648 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1649 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1650 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1651 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1652 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1653 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1654 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1655 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1656 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1657 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1658 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1659 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1660 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1661 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1662 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1663 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1664 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1665 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1666 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1667 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1668 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1669 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1670 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1671 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1672 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1673 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1674 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1675 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1676 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1677 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1678 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1679 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1680 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1681 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1682 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1683 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1684 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1685 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1686 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1687 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1688 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1689 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1690 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1691 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1692 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1693 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1694 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1695 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1696 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1697 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1698 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1699 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1700 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1701 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1702 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1703 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1704 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1705 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1706 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1707 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1708 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1709 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1710 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1711 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1712 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1713 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1714 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1715 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1716 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1717 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1718 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1719 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1720 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1721 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1722 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1723 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1724 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1725 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1726 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1727 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1728 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1729 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1730 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1731 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1732 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1733 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1734 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1735 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1736 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1737 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1738 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1739 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1740 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1741 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1742 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1743 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1744 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1745 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1746 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1747 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1748 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1749 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1750 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1751 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1752 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1753 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1754 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1755 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1756 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1757 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1758 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1759 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1760 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1761 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1762 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1763 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1764 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1765 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1766 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1767 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1768 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1769 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1770 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1771 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1772 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1773 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1774 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1775 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1776 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1777 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1778 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1779 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1780 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1781 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1782 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1783 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1784 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1785 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1786 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1787 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1788 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1789 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1790 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1791 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1792 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1793 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1794 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1795 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1796 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1797 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1798 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1799 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1800 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1801 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1802 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1803 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1804 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1805 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1806 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1807 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1808 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1809 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1810 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1811 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1812 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1813 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1814 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1815 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1816 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1817 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1818 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1819 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1820 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1821 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1822 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1823 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1824 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1825 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1826 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1827 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1828 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1829 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1830 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1831 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1832 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1833 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1834 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1835 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1836 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1837 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1838 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1839 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1840 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1841 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1842 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1843 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1844 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1845 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1846 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1847 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1848 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1849 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1850 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1851 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1852 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1853 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1854 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1855 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1856 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1857 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1858 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1859 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1860 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1861 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1862 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1863 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1864 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1865 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1866 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1867 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1868 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1869 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1870 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1871 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1872 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1873 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1874 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1875 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1876 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1877 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1878 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1879 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1880 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1881 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1882 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1883 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1884 outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1885 OutputP V_da2_P outd_stage3_0/outd_stage2_0/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1886 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1887 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1888 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1889 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1890 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1891 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1892 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1893 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1894 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1895 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1896 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1897 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1898 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1899 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1900 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1901 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1902 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1903 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1904 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1905 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1906 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1907 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1908 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1909 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1910 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1911 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1912 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1913 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1914 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1915 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1916 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1917 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1918 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1919 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1920 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1921 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1922 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1923 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1924 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1925 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1926 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1927 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1928 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1929 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1930 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1931 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1932 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1933 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1934 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1935 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1936 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1937 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1938 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1939 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1940 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1941 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1942 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1943 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1944 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1945 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1946 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1947 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1948 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1949 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1950 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1951 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1952 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1953 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1954 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1955 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1956 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1957 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1958 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1959 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1960 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1961 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1962 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1963 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1964 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1965 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1966 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1967 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1968 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1969 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1970 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1971 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1972 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1973 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1974 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1975 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1976 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1977 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1978 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1979 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1980 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1981 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1982 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1983 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1984 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1985 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1986 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1987 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1988 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1989 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1990 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1991 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1992 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1993 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1994 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1995 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1996 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1997 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1998 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1999 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2000 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2001 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2002 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2003 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2004 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2005 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2006 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2007 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2008 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2009 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2010 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2011 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2012 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2013 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2014 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2015 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2016 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2017 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2018 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2019 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2020 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2021 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2022 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2023 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2024 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2025 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2026 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2027 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2028 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2029 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2030 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2031 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2032 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2033 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2034 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2035 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2036 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2037 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2038 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2039 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2040 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2041 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2042 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2043 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2044 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2045 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2046 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2047 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2048 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2049 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2050 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2051 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2052 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2053 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2054 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2055 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2056 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2057 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2058 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2059 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2060 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2061 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2062 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2063 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2064 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2065 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2066 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2067 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2068 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2069 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2070 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2071 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2072 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2073 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2074 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2075 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2076 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2077 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2078 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2079 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2080 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2081 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2082 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2083 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2084 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2085 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2086 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2087 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2088 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2089 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2090 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2091 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2092 VN V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2093 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2094 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2095 VN V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2096 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2097 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2098 outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2099 OutputN V_da2_N outd_stage3_0/outd_stage2_0/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2100 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2101 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2102 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2103 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2104 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2105 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2106 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2107 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2108 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2109 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2110 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2111 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2112 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2113 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2114 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2115 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2116 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2117 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2118 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2119 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2120 VN V_da2_P OutputP outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2121 OutputP V_da2_P VN outd_stage3_0/outd_stage2_0/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2122 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2123 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2124 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2125 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2126 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2127 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2128 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2129 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2130 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2131 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2132 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2133 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2134 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2135 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2136 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2137 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2138 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2139 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2140 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2141 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2142 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2143 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2144 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2145 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2146 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2147 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2148 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2149 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2150 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2151 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2152 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2153 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2154 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2155 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2156 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2157 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2158 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2159 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2160 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2161 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2162 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2163 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2164 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2165 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2166 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2167 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2168 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2169 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2170 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2171 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2172 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2173 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2174 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2175 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2176 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2177 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2178 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2179 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2180 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2181 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2182 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2183 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2184 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2185 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2186 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2187 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2188 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2189 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2190 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2191 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2192 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2193 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2194 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2195 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2196 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2197 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2198 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2199 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2200 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2201 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2202 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2203 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2204 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2205 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2206 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2207 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2208 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2209 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2210 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2211 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2212 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2213 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2214 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2215 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2216 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2217 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2218 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2219 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2220 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2221 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2222 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2223 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2224 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2225 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2226 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2227 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2228 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2229 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2230 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2231 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2232 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2233 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2234 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2235 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2236 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2237 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2238 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2239 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2240 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2241 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2242 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2243 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2244 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2245 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2246 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2247 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2248 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2249 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2250 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2251 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2252 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2253 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2254 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2255 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2256 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2257 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2258 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2259 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2260 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2261 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2262 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2263 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2264 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2265 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2266 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2267 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2268 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2269 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2270 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2271 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2272 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2273 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2274 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2275 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2276 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2277 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2278 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2279 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2280 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2281 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2282 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2283 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2284 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2285 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2286 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2287 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2288 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2289 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2290 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2291 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2292 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2293 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2294 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2295 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2296 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2297 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2298 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2299 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2300 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2301 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2302 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2303 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2304 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2305 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2306 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2307 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2308 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2309 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2310 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2311 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2312 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2313 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2314 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2315 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2316 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2317 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2318 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2319 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2320 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2321 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2322 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2323 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2324 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2325 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2326 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2327 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2328 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2329 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2330 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2331 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2332 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2333 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2334 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2335 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2336 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2337 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2338 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2339 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2340 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2341 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2342 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2343 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2344 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2345 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2346 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2347 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2348 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2349 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2350 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2351 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2352 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2353 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2354 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2355 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2356 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2357 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2358 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2359 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2360 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2361 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2362 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2363 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2364 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2365 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2366 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2367 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2368 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2369 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2370 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2371 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2372 outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2373 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2374 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2375 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2376 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2377 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2378 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2379 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2380 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2381 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2382 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2383 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2384 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2385 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2386 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2387 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2388 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2389 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2390 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2391 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2392 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2393 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2394 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2395 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2396 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2397 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2398 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2399 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2400 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2401 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2402 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2403 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2404 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2405 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2406 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2407 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2408 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2409 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2410 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2411 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2412 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2413 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2414 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2415 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2416 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2417 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2418 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2419 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2420 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2421 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2422 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2423 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2424 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2425 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2426 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2427 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2428 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2429 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2430 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2431 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2432 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2433 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2434 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2435 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2436 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2437 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2438 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2439 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2440 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2441 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2442 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2443 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2444 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2445 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2446 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2447 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2448 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2449 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2450 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2451 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2452 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2453 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2454 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2455 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2456 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2457 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2458 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2459 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2460 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2461 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2462 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2463 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2464 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2465 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2466 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2467 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2468 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2469 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2470 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2471 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2472 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2473 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2474 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2475 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2476 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2477 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2478 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2479 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2480 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2481 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2482 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2483 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2484 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2485 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2486 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2487 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2488 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2489 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2490 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2491 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2492 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2493 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2494 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2495 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2496 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2497 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2498 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2499 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2500 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2501 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2502 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2503 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2504 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2505 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2506 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2507 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2508 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2509 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2510 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2511 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2512 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2513 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2514 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2515 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2516 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2517 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2518 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2519 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2520 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2521 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2522 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2523 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2524 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2525 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2526 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2527 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2528 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2529 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2530 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2531 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2532 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2533 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2534 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2535 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2536 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2537 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2538 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2539 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2540 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2541 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2542 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2543 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2544 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2545 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2546 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2547 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2548 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2549 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2550 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2551 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2552 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2553 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2554 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2555 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2556 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2557 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2558 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2559 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2560 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2561 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2562 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2563 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2564 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2565 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2566 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2567 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2568 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2569 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2570 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2571 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2572 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2573 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2574 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2575 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2576 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2577 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2578 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2579 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2580 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2581 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2582 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2583 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2584 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2585 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2586 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2587 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2588 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2589 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2590 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2591 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2592 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2593 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2594 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2595 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2596 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2597 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2598 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2599 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2600 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2601 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2602 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2603 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2604 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2605 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2606 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2607 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2608 outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2609 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2610 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2611 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2612 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2613 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2614 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2615 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2616 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2617 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2618 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2619 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2620 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2621 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2622 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2623 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2624 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2625 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2626 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2627 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2628 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2629 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2630 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2631 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2632 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2633 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2634 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2635 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2636 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2637 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2638 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2639 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2640 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2641 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2642 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2643 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2644 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2645 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2646 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2647 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2648 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2649 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2650 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2651 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2652 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2653 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2654 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2655 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2656 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2657 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2658 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2659 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2660 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2661 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2662 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2663 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2664 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2665 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2666 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2667 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2668 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2669 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2670 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2671 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2672 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2673 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2674 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2675 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2676 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2677 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2678 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2679 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2680 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2681 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2682 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2683 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2684 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2685 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2686 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2687 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2688 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2689 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2690 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2691 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2692 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2693 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2694 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2695 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2696 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2697 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2698 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2699 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2700 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2701 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2702 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2703 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2704 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2705 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2706 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2707 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2708 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2709 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2710 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2711 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2712 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2713 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2714 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2715 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2716 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2717 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2718 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2719 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2720 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2721 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2722 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2723 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2724 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2725 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2726 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2727 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2728 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2729 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2730 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2731 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2732 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2733 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2734 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2735 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2736 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2737 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2738 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2739 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2740 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2741 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2742 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2743 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2744 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2745 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2746 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2747 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2748 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2749 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2750 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2751 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2752 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2753 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2754 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2755 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2756 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2757 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2758 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2759 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2760 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2761 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2762 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2763 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2764 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2765 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2766 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2767 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2768 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2769 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2770 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2771 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2772 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2773 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2774 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2775 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2776 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2777 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2778 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2779 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2780 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2781 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2782 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2783 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2784 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2785 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2786 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2787 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2788 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2789 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2790 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2791 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2792 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2793 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2794 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2795 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2796 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2797 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2798 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2799 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2800 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2801 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2802 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2803 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2804 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2805 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2806 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2807 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2808 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2809 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2810 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2811 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2812 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2813 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2814 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2815 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2816 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2817 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2818 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2819 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2820 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2821 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2822 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2823 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2824 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2825 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2826 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2827 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2828 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2829 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2830 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2831 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2832 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2833 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2834 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2835 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2836 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2837 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2838 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2839 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2840 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2841 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2842 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2843 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2844 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2845 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2846 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2847 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2848 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2849 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2850 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2851 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2852 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2853 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2854 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2855 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2856 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2857 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2858 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2859 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2860 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2861 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2862 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2863 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2864 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2865 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2866 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2867 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2868 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2869 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2870 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2871 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2872 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2873 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2874 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2875 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2876 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2877 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2878 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2879 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2880 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2881 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2882 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2883 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2884 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2885 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2886 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2887 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2888 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2889 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2890 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2891 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2892 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2893 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2894 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2895 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2896 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2897 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2898 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2899 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2900 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2901 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2902 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2903 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2904 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2905 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2906 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2907 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2908 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2909 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2910 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2911 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2912 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2913 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2914 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2915 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2916 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2917 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2918 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2919 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2920 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2921 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2922 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2923 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2924 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2925 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2926 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2927 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2928 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2929 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2930 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2931 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2932 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2933 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2934 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2935 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2936 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2937 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2938 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2939 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2940 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2941 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2942 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2943 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2944 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2945 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2946 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2947 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2948 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2949 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2950 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2951 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2952 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2953 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2954 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2955 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2956 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2957 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2958 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2959 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2960 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2961 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2962 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2963 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2964 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2965 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2966 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2967 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2968 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2969 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2970 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2971 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2972 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2973 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2974 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2975 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2976 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2977 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2978 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2979 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2980 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2981 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2982 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2983 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2984 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2985 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2986 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2987 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2988 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2989 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2990 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2991 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2992 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2993 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2994 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2995 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2996 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2997 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2998 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2999 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3000 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3001 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3002 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3003 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3004 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3005 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3006 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3007 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3008 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3009 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3010 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3011 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3012 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3013 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3014 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3015 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3016 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3017 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3018 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3019 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3020 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3021 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3022 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3023 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3024 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3025 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3026 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3027 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3028 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3029 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3030 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3031 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3032 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3033 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3034 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3035 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3036 outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3037 OutputP V_da2_P outd_stage3_0/outd_stage2_1/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3038 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3039 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3040 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3041 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3042 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3043 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3044 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3045 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3046 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3047 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3048 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3049 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3050 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3051 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3052 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3053 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3054 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3055 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3056 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3057 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3058 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3059 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3060 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3061 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3062 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3063 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3064 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3065 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3066 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3067 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3068 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3069 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3070 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3071 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3072 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3073 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3074 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3075 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3076 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3077 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3078 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3079 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3080 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3081 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3082 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3083 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3084 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3085 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3086 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3087 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3088 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3089 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3090 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3091 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3092 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3093 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3094 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3095 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3096 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3097 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3098 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3099 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3100 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3101 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3102 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3103 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3104 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3105 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3106 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3107 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3108 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3109 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3110 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3111 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3112 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3113 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3114 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3115 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3116 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3117 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3118 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3119 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3120 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3121 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3122 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3123 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3124 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3125 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3126 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3127 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3128 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3129 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3130 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3131 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3132 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3133 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3134 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3135 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3136 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3137 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3138 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3139 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3140 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3141 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3142 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3143 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3144 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3145 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3146 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3147 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3148 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3149 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3150 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3151 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3152 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3153 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3154 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3155 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3156 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3157 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3158 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3159 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3160 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3161 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3162 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3163 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3164 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3165 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3166 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3167 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3168 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3169 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3170 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3171 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3172 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3173 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3174 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3175 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3176 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3177 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3178 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3179 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3180 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3181 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3182 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3183 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3184 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3185 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3186 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3187 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3188 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3189 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3190 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3191 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3192 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3193 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3194 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3195 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3196 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3197 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3198 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3199 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3200 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3201 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3202 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3203 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3204 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3205 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3206 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3207 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3208 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3209 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3210 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3211 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3212 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3213 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3214 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3215 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3216 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3217 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3218 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3219 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3220 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3221 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3222 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3223 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3224 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3225 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3226 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3227 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3228 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3229 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3230 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3231 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3232 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3233 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3234 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3235 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3236 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3237 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3238 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3239 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3240 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3241 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3242 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3243 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3244 VN V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3245 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3246 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3247 VN V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3248 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3249 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3250 outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3251 OutputN V_da2_N outd_stage3_0/outd_stage2_1/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3252 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3253 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3254 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3255 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3256 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3257 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3258 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3259 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3260 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3261 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3262 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3263 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3264 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3265 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3266 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3267 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3268 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3269 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3270 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3271 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3272 VN V_da2_P OutputP outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3273 OutputP V_da2_P VN outd_stage3_0/outd_stage2_1/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3274 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3275 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3276 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3277 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3278 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3279 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3280 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3281 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3282 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3283 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3284 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3285 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3286 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3287 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3288 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3289 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3290 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3291 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3292 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3293 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3294 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3295 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3296 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3297 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3298 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3299 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3300 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3301 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3302 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3303 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3304 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3305 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3306 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3307 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3308 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3309 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3310 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3311 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3312 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3313 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3314 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3315 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3316 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3317 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3318 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3319 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3320 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3321 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3322 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3323 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3324 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3325 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3326 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3327 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3328 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3329 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3330 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3331 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3332 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3333 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3334 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3335 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3336 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3337 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3338 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3339 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3340 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3341 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3342 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3343 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3344 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3345 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3346 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3347 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3348 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3349 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3350 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3351 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3352 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3353 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3354 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3355 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3356 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3357 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3358 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3359 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3360 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3361 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3362 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3363 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3364 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3365 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3366 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3367 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3368 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3369 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3370 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3371 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3372 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3373 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3374 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3375 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3376 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3377 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3378 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3379 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3380 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3381 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3382 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3383 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3384 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3385 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3386 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3387 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3388 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3389 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3390 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3391 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3392 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3393 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3394 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3395 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3396 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3397 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3398 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3399 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3400 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3401 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3402 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3403 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3404 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3405 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3406 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3407 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3408 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3409 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3410 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3411 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3412 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3413 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3414 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3415 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3416 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3417 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3418 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3419 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3420 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3421 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3422 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3423 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3424 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3425 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3426 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3427 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3428 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3429 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3430 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3431 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3432 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3433 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3434 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3435 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3436 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3437 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3438 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3439 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3440 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3441 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3442 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3443 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3444 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3445 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3446 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3447 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3448 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3449 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3450 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3451 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3452 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3453 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3454 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3455 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3456 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3457 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3458 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3459 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3460 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3461 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3462 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3463 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3464 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3465 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3466 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3467 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3468 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3469 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3470 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3471 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3472 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3473 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3474 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3475 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3476 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3477 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3478 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3479 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3480 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3481 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3482 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3483 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3484 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3485 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3486 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3487 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3488 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3489 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3490 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3491 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3492 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3493 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3494 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3495 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3496 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3497 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3498 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3499 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3500 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3501 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3502 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3503 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3504 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3505 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3506 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3507 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3508 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3509 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3510 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3511 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3512 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3513 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3514 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3515 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3516 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3517 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3518 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3519 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3520 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3521 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3522 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3523 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3524 outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3525 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3526 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3527 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3528 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3529 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3530 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3531 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3532 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3533 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3534 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3535 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3536 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3537 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3538 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3539 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3540 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3541 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3542 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3543 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3544 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3545 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3546 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3547 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3548 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3549 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3550 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3551 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3552 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3553 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3554 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3555 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3556 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3557 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3558 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3559 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3560 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3561 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3562 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3563 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3564 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3565 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3566 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3567 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3568 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3569 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3570 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3571 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3572 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3573 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3574 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3575 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3576 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3577 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3578 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3579 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3580 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3581 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3582 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3583 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3584 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3585 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3586 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3587 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3588 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3589 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3590 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3591 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3592 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3593 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3594 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3595 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3596 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3597 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3598 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3599 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3600 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3601 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3602 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3603 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3604 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3605 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3606 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3607 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3608 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3609 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3610 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3611 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3612 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3613 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3614 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3615 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3616 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3617 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3618 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3619 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3620 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3621 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3622 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3623 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3624 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3625 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3626 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3627 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3628 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3629 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3630 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3631 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3632 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3633 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3634 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3635 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3636 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3637 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3638 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3639 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3640 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3641 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3642 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3643 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3644 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3645 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3646 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3647 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3648 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3649 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3650 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3651 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3652 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3653 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3654 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3655 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3656 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3657 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3658 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3659 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3660 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3661 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3662 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3663 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3664 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3665 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3666 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3667 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3668 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3669 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3670 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3671 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3672 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3673 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3674 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3675 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3676 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3677 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3678 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3679 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3680 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3681 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3682 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3683 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3684 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3685 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3686 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3687 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3688 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3689 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3690 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3691 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3692 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3693 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3694 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3695 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3696 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3697 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3698 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3699 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3700 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3701 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3702 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3703 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3704 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3705 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3706 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3707 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3708 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3709 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3710 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3711 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3712 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3713 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3714 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3715 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3716 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3717 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3718 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3719 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3720 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3721 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3722 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3723 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3724 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3725 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3726 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3727 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3728 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3729 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3730 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3731 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3732 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3733 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3734 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3735 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3736 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3737 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3738 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3739 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3740 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3741 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3742 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3743 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3744 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3745 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3746 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3747 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3748 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3749 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3750 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3751 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3752 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3753 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3754 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3755 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3756 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3757 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3758 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3759 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3760 outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3761 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3762 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3763 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3764 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3765 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3766 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3767 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3768 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3769 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3770 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3771 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3772 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3773 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3774 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3775 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3776 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3777 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3778 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3779 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3780 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3781 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3782 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3783 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3784 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3785 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3786 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3787 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3788 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3789 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3790 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3791 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3792 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3793 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3794 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3795 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3796 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3797 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3798 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3799 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3800 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3801 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3802 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3803 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3804 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3805 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3806 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3807 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3808 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3809 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3810 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3811 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3812 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3813 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3814 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3815 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3816 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3817 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3818 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3819 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3820 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3821 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3822 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3823 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3824 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3825 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3826 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3827 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3828 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3829 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3830 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3831 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3832 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3833 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3834 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3835 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3836 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3837 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3838 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3839 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3840 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3841 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3842 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3843 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3844 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3845 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3846 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3847 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3848 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3849 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3850 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3851 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3852 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3853 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3854 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3855 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3856 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3857 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3858 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3859 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3860 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3861 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3862 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3863 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3864 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3865 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3866 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3867 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3868 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3869 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3870 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3871 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3872 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3873 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3874 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3875 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3876 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3877 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3878 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3879 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3880 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3881 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3882 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3883 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3884 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3885 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3886 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3887 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3888 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3889 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3890 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3891 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3892 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3893 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3894 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3895 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3896 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3897 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3898 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3899 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3900 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3901 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3902 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3903 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3904 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3905 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3906 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3907 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3908 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3909 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3910 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3911 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3912 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3913 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3914 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3915 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3916 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3917 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3918 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3919 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3920 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3921 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3922 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3923 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3924 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3925 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3926 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3927 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3928 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3929 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3930 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3931 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3932 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3933 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3934 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3935 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3936 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3937 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3938 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3939 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3940 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3941 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3942 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3943 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3944 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3945 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3946 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3947 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3948 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3949 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3950 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3951 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3952 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3953 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3954 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3955 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3956 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3957 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3958 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3959 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3960 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3961 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3962 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3963 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3964 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3965 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3966 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3967 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3968 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3969 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3970 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3971 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3972 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3973 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3974 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3975 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3976 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3977 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3978 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3979 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3980 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3981 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3982 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3983 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3984 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3985 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3986 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3987 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3988 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3989 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3990 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3991 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3992 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3993 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3994 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3995 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3996 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3997 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3998 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3999 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4000 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4001 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4002 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4003 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4004 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4005 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4006 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4007 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4008 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4009 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4010 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4011 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4012 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4013 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4014 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4015 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4016 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4017 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4018 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4019 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4020 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4021 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4022 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4023 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4024 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4025 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4026 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4027 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4028 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4029 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4030 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4031 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4032 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4033 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4034 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4035 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4036 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4037 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4038 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4039 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4040 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4041 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4042 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4043 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4044 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4045 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4046 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4047 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4048 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4049 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4050 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4051 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4052 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4053 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4054 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4055 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4056 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4057 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4058 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4059 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4060 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4061 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4062 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4063 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4064 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4065 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4066 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4067 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4068 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4069 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4070 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4071 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4072 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4073 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4074 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4075 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4076 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4077 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4078 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4079 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4080 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4081 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4082 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4083 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4084 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4085 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4086 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4087 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4088 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4089 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4090 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4091 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4092 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4093 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4094 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4095 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4096 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4097 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4098 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4099 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4100 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4101 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4102 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4103 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4104 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4105 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4106 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4107 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4108 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4109 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4110 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4111 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4112 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4113 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4114 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4115 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4116 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4117 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4118 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4119 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4120 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4121 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4122 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4123 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4124 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4125 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4126 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4127 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4128 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4129 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4130 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4131 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4132 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4133 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4134 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4135 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4136 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4137 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4138 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4139 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4140 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4141 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4142 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4143 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4144 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4145 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4146 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4147 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4148 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4149 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4150 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4151 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4152 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4153 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4154 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4155 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4156 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4157 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4158 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4159 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4160 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4161 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4162 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4163 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4164 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4165 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4166 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4167 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4168 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4169 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4170 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4171 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4172 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4173 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4174 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4175 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4176 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4177 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4178 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4179 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4180 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4181 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4182 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4183 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4184 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4185 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4186 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4187 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4188 outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4189 OutputP V_da2_P outd_stage3_0/outd_stage2_2/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4190 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4191 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4192 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4193 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4194 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4195 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4196 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4197 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4198 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4199 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4200 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4201 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4202 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4203 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4204 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4205 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4206 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4207 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4208 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4209 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4210 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4211 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4212 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4213 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4214 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4215 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4216 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4217 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4218 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4219 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4220 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4221 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4222 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4223 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4224 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4225 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4226 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4227 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4228 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4229 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4230 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4231 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4232 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4233 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4234 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4235 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4236 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4237 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4238 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4239 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4240 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4241 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4242 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4243 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4244 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4245 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4246 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4247 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4248 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4249 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4250 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4251 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4252 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4253 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4254 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4255 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4256 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4257 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4258 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4259 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4260 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4261 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4262 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4263 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4264 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4265 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4266 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4267 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4268 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4269 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4270 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4271 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4272 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4273 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4274 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4275 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4276 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4277 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4278 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4279 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4280 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4281 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4282 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4283 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4284 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4285 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4286 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4287 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4288 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4289 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4290 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4291 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4292 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4293 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4294 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4295 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4296 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4297 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4298 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4299 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4300 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4301 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4302 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4303 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4304 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4305 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4306 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4307 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4308 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4309 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4310 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4311 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4312 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4313 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4314 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4315 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4316 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4317 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4318 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4319 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4320 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4321 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4322 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4323 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4324 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4325 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4326 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4327 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4328 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4329 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4330 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4331 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4332 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4333 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4334 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4335 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4336 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4337 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4338 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4339 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4340 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4341 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4342 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4343 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4344 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4345 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4346 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4347 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4348 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4349 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4350 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4351 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4352 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4353 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4354 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4355 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4356 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4357 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4358 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4359 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4360 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4361 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4362 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4363 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4364 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4365 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4366 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4367 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4368 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4369 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4370 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4371 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4372 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4373 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4374 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4375 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4376 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4377 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4378 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4379 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4380 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4381 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4382 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4383 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4384 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4385 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4386 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4387 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4388 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4389 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4390 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4391 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4392 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4393 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4394 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4395 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4396 VN V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4397 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4398 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4399 VN V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4400 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4401 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4402 outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4403 OutputN V_da2_N outd_stage3_0/outd_stage2_2/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4404 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4405 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4406 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4407 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4408 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4409 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4410 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4411 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4412 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4413 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4414 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4415 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4416 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4417 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4418 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4419 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4420 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4421 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4422 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4423 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4424 VN V_da2_P OutputP outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4425 OutputP V_da2_P VN outd_stage3_0/outd_stage2_2/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4426 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4427 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4428 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4429 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4430 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4431 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4432 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4433 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4434 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4435 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4436 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4437 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4438 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4439 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4440 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4441 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4442 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4443 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4444 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4445 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4446 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4447 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4448 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4449 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4450 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4451 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4452 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4453 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4454 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4455 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4456 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4457 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4458 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4459 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4460 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4461 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4462 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4463 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4464 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4465 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4466 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4467 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4468 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4469 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4470 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4471 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4472 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4473 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4474 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4475 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4476 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4477 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4478 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4479 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4480 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4481 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4482 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4483 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4484 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4485 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4486 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4487 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4488 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4489 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4490 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4491 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4492 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4493 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4494 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4495 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4496 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4497 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4498 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4499 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4500 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4501 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4502 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4503 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4504 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4505 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4506 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4507 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4508 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4509 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4510 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4511 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4512 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4513 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4514 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4515 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4516 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4517 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4518 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4519 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4520 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4521 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4522 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4523 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4524 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4525 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4526 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4527 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4528 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4529 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4530 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4531 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4532 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4533 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4534 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4535 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4536 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4537 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4538 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4539 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4540 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4541 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4542 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4543 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4544 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4545 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4546 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4547 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4548 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4549 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4550 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4551 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4552 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4553 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4554 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4555 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4556 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4557 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4558 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4559 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4560 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4561 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4562 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4563 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4564 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4565 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4566 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4567 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4568 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4569 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4570 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4571 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4572 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4573 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4574 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4575 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4576 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4577 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4578 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4579 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4580 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4581 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4582 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4583 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4584 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4585 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4586 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4587 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4588 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4589 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4590 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4591 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4592 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4593 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4594 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4595 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4596 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4597 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4598 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4599 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4600 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4601 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4602 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4603 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4604 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4605 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4606 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4607 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4608 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4609 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4610 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4611 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4612 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4613 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4614 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4615 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4616 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4617 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4618 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4619 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4620 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4621 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4622 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4623 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4624 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4625 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4626 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4627 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4628 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4629 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4630 VP OutputP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4631 VP OutputN VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4632 OutputN VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4633 OutputP VP VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4634 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4635 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4636 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4637 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4638 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4639 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4640 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4641 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4642 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4643 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4644 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4645 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4646 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4647 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4648 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4649 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4650 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4651 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4652 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4653 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4654 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4655 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4656 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4657 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4658 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4659 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4660 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4661 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4662 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4663 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4664 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4665 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4666 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4667 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4668 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4669 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4670 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4671 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4672 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4673 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4674 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4675 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4676 outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4677 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_0/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_0/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4678 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4679 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4680 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4681 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4682 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4683 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4684 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4685 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4686 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4687 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4688 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4689 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4690 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4691 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4692 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4693 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4694 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4695 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4696 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4697 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4698 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4699 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4700 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4701 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4702 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4703 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4704 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4705 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4706 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4707 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4708 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4709 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4710 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4711 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4712 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4713 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4714 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4715 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4716 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4717 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4718 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4719 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4720 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4721 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4722 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4723 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4724 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4725 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4726 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4727 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4728 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4729 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4730 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4731 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4732 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4733 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4734 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4735 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4736 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4737 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4738 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4739 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4740 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4741 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4742 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4743 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4744 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4745 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4746 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4747 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4748 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4749 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4750 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4751 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4752 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4753 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4754 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4755 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4756 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4757 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4758 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4759 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4760 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4761 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4762 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4763 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4764 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4765 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4766 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4767 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4768 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4769 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4770 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4771 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4772 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4773 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4774 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4775 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4776 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4777 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4778 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4779 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4780 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4781 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4782 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4783 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4784 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4785 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4786 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4787 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4788 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4789 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4790 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4791 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4792 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4793 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4794 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4795 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4796 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4797 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4798 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4799 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4800 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4801 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4802 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4803 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4804 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4805 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4806 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4807 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4808 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4809 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4810 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4811 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4812 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4813 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4814 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4815 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4816 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4817 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4818 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4819 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4820 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4821 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4822 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4823 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4824 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4825 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4826 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4827 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4828 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4829 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4830 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4831 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4832 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4833 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4834 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4835 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4836 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4837 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4838 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4839 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4840 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4841 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4842 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4843 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4844 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4845 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4846 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4847 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4848 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4849 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4850 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4851 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4852 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4853 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4854 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4855 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4856 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4857 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4858 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4859 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4860 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4861 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4862 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4863 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4864 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4865 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4866 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4867 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4868 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4869 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4870 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4871 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4872 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4873 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4874 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4875 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4876 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4877 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4878 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4879 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4880 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4881 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4882 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4883 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4884 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4885 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4886 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4887 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4888 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4889 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4890 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4891 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4892 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4893 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4894 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4895 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4896 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4897 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4898 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4899 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4900 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4901 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4902 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4903 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4904 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4905 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4906 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4907 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4908 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4909 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4910 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4911 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4912 outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4913 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_1/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_1/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4914 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4915 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4916 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4917 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4918 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4919 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4920 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4921 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4922 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4923 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4924 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4925 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4926 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4927 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4928 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4929 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4930 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4931 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4932 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4933 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4934 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4935 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4936 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4937 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4938 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4939 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4940 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4941 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4942 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4943 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4944 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4945 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4946 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4947 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4948 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4949 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4950 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4951 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4952 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4953 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4954 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4955 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4956 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4957 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4958 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4959 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4960 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4961 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4962 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4963 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4964 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4965 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4966 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4967 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4968 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4969 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4970 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4971 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4972 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4973 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4974 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4975 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4976 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4977 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4978 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4979 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4980 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4981 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4982 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4983 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4984 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4985 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4986 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4987 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4988 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4989 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4990 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4991 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4992 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4993 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4994 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4995 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4996 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4997 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4998 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4999 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5000 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5001 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5002 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5003 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5004 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5005 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5006 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5007 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5008 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5009 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5010 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5011 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5012 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5013 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5014 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5015 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5016 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5017 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5018 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5019 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5020 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5021 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5022 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5023 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5024 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5025 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5026 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5027 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5028 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5029 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5030 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5031 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5032 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5033 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5034 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5035 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5036 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5037 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5038 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5039 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5040 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5041 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5042 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5043 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5044 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5045 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5046 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5047 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5048 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5049 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5050 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5051 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5052 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5053 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5054 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5055 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5056 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5057 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5058 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5059 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5060 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5061 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5062 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5063 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5064 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5065 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5066 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5067 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5068 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5069 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5070 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5071 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5072 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5073 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5074 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5075 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5076 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5077 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5078 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5079 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5080 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5081 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5082 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5083 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5084 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5085 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5086 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5087 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5088 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5089 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5090 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5091 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5092 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5093 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5094 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5095 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5096 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5097 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5098 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5099 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5100 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5101 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5102 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5103 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5104 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5105 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5106 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5107 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5108 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5109 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5110 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5111 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5112 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5113 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5114 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5115 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5116 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5117 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5118 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5119 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5120 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5121 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5122 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5123 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5124 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5125 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5126 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5127 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5128 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5129 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5130 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5131 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5132 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5133 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5134 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5135 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5136 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5137 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5138 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5139 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5140 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5141 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5142 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5143 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5144 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5145 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5146 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5147 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5148 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5149 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5150 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5151 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5152 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5153 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5154 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5155 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5156 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5157 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5158 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5159 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5160 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5161 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5162 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5163 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5164 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5165 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5166 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5167 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5168 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5169 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5170 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5171 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5172 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5173 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5174 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5175 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5176 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5177 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5178 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5179 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5180 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5181 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5182 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5183 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5184 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5185 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5186 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5187 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5188 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5189 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5190 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5191 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5192 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5193 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5194 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5195 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5196 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5197 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5198 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5199 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5200 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5201 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5202 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5203 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5204 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5205 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5206 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5207 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5208 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5209 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5210 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5211 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5212 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5213 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5214 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5215 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5216 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5217 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5218 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5219 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5220 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5221 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5222 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5223 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5224 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5225 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5226 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5227 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5228 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5229 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5230 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5231 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5232 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5233 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5234 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5235 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5236 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5237 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5238 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5239 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5240 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5241 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5242 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5243 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5244 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5245 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5246 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5247 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5248 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5249 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5250 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5251 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5252 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5253 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5254 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5255 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5256 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5257 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5258 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5259 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5260 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5261 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5262 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5263 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5264 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5265 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5266 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5267 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5268 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5269 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5270 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5271 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5272 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5273 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5274 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5275 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5276 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5277 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5278 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5279 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5280 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5281 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5282 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5283 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5284 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5285 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5286 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5287 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5288 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5289 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5290 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5291 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5292 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5293 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5294 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5295 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5296 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5297 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5298 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5299 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5300 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5301 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5302 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5303 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5304 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5305 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5306 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5307 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5308 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5309 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5310 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5311 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5312 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5313 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5314 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5315 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5316 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5317 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5318 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5319 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5320 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5321 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5322 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5323 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5324 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5325 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5326 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5327 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5328 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5329 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5330 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5331 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5332 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5333 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5334 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5335 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5336 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5337 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5338 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5339 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5340 outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5341 OutputP V_da2_P outd_stage3_0/outd_stage2_3/outd_diffamp_2/m1_2468_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_2/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5342 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5343 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5344 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5345 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5346 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5347 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5348 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5349 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5350 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5351 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5352 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5353 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5354 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5355 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5356 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5357 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5358 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5359 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5360 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5361 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5362 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5363 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5364 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5365 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5366 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5367 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5368 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5369 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5370 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5371 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5372 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5373 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5374 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5375 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5376 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5377 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5378 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5379 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5380 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5381 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5382 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5383 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5384 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5385 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5386 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5387 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5388 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5389 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5390 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5391 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5392 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5393 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5394 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5395 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5396 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5397 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5398 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5399 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5400 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5401 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5402 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5403 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5404 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5405 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5406 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5407 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5408 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5409 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5410 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5411 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5412 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5413 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5414 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5415 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5416 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5417 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5418 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5419 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5420 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5421 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5422 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5423 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5424 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5425 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5426 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5427 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5428 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5429 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5430 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5431 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5432 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5433 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5434 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5435 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5436 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5437 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5438 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5439 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5440 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5441 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5442 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5443 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5444 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5445 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5446 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5447 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5448 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5449 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5450 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5451 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5452 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5453 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5454 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5455 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5456 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5457 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5458 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5459 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5460 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5461 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5462 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5463 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5464 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5465 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5466 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5467 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5468 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5469 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5470 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5471 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5472 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5473 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5474 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5475 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5476 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5477 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5478 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5479 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5480 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5481 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5482 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5483 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5484 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5485 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5486 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5487 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5488 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5489 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5490 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5491 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5492 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5493 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5494 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5495 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5496 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5497 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5498 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5499 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5500 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5501 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5502 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5503 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5504 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5505 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5506 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5507 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5508 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5509 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5510 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5511 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5512 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5513 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5514 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5515 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5516 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5517 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5518 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5519 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5520 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5521 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5522 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5523 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5524 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5525 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5526 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5527 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5528 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5529 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5530 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5531 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5532 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5533 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5534 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5535 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5536 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5537 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5538 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5539 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5540 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5541 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5542 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5543 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5544 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5545 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5546 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5547 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5548 VN V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5549 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5550 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5551 VN V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5552 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5553 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5554 outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# V_da2_N OutputN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5555 OutputN V_da2_N outd_stage3_0/outd_stage2_3/outd_diffamp_3/m1_994_8758# outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5556 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5557 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5558 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5559 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5560 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5561 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5562 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5563 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5564 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5565 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5566 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5567 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5568 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5569 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5570 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5571 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5572 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5573 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5574 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5575 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5576 VN V_da2_P OutputP outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5577 OutputP V_da2_P VN outd_stage3_0/outd_stage2_3/outd_diffamp_3/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5578 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5579 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5580 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5581 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5582 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5583 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5584 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5585 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5586 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5587 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5588 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5589 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5590 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5591 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5592 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5593 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5594 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5595 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5596 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5597 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5598 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5599 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5600 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5601 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5602 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5603 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5604 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5605 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5606 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5607 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5608 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5609 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5610 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5611 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5612 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5613 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5614 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5615 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5616 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5617 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5618 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5619 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5620 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5621 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5622 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5623 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5624 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5625 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5626 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5627 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5628 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5629 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5630 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5631 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5632 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5633 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5634 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5635 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5636 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5637 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5638 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5639 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5640 VM14D I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5641 outd_stage3_0/m2_41490_8160# I_Bias VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5642 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5643 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5644 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5645 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5646 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5647 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5648 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5649 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5650 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5651 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5652 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5653 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5654 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5655 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5656 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5657 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5658 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5659 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5660 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5661 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5662 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5663 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5664 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5665 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5666 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5667 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5668 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5669 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5670 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5671 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5672 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5673 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5674 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5675 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5676 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5677 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5678 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5679 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5680 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5681 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5682 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5683 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5684 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5685 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5686 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5687 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5688 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5689 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5690 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5691 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5692 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5693 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5694 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5695 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5696 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5697 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5698 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5699 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5700 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5701 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5702 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5703 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5704 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5705 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5706 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5707 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5708 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5709 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5710 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5711 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5712 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5713 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5714 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5715 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5716 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5717 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5718 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5719 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5720 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5721 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5722 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5723 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5724 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5725 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5726 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5727 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5728 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5729 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5730 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5731 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5732 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5733 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5734 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5735 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5736 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5737 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5738 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5739 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5740 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5741 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5742 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5743 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5744 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5745 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5746 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5747 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5748 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5749 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5750 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5751 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5752 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5753 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5754 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5755 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5756 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5757 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5758 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5759 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5760 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5761 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5762 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5763 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5764 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5765 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5766 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5767 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5768 VN I_Bias outd_stage3_0/m2_41490_8160# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5769 outd_stage3_0/m2_41490_8160# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5770 I_Bias I_Bias m1_n19890_7120# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5771 m1_n19890_7120# I_Bias I_Bias VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5772 InputRef VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5773 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5774 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5775 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5776 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5777 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5778 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5779 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5780 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5781 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5782 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5783 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5784 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5785 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5786 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5787 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5788 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5789 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5790 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5791 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5792 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5793 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5794 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5795 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5796 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5797 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5798 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5799 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5800 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5801 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5802 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5803 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5804 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5805 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5806 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5807 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5808 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5809 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5810 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5811 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5812 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5813 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5814 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5815 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5816 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5817 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5818 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5819 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5820 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5821 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5822 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5823 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5824 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5825 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5826 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5827 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5828 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5829 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5830 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5831 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5832 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5833 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5834 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5835 outd_stage1_0/isource_out I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5836 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias outd_stage1_0/isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5837 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5838 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5839 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5840 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5841 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5842 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5843 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5844 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5845 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5846 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5847 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5848 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5849 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5850 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5851 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5852 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5853 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5854 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5855 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5856 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5857 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5858 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5859 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5860 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5861 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5862 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5863 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5864 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5865 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5866 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5867 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5868 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5869 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5870 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5871 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5872 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5873 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5874 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5875 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5876 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5877 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5878 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5879 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5880 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5881 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5882 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5883 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5884 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5885 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5886 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5887 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5888 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5889 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5890 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5891 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5892 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5893 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5894 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5895 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5896 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5897 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5898 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5899 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5900 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5901 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5902 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5903 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5904 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5905 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5906 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5907 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5908 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5909 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5910 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5911 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5912 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5913 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5914 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5915 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5916 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5917 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5918 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5919 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5920 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5921 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5922 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5923 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5924 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5925 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5926 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5927 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5928 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5929 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5930 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5931 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5932 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5933 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5934 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5935 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5936 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5937 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5938 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5939 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5940 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5941 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5942 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5943 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5944 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5945 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5946 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5947 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5948 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5949 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5950 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5951 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5952 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5953 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5954 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5955 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5956 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5957 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5958 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5959 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5960 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5961 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5962 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5963 VN I_Bias outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5964 outd_stage1_0/outd_cmirror_64t_0/m1_220_5610# I_Bias VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5965 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5966 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5967 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5968 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5969 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5970 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5971 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5972 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5973 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5974 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5975 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5976 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5977 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5978 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5979 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5980 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5981 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5982 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5983 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5984 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5985 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5986 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5987 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5988 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5989 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5990 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5991 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5992 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5993 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5994 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5995 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5996 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5997 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5998 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5999 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6000 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6001 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6002 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6003 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6004 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6005 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6006 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6007 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6008 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6009 V_da1_P VP VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6010 V_da1_P VP VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6011 V_da1_P VP VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6012 V_da1_P VP VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6013 V_da1_N VP VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6014 V_da1_N VP VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6015 V_da1_N VP VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6016 V_da1_N VP VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X6017 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6018 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6019 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6020 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6021 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6022 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
