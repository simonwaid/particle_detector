magic
tech sky130A
magscale 1 2
timestamp 1645790779
<< error_p >>
rect -1181 581 -1123 587
rect -989 581 -931 587
rect -797 581 -739 587
rect -605 581 -547 587
rect -413 581 -355 587
rect -221 581 -163 587
rect -29 581 29 587
rect 163 581 221 587
rect 355 581 413 587
rect 547 581 605 587
rect 739 581 797 587
rect 931 581 989 587
rect 1123 581 1181 587
rect -1181 547 -1169 581
rect -989 547 -977 581
rect -797 547 -785 581
rect -605 547 -593 581
rect -413 547 -401 581
rect -221 547 -209 581
rect -29 547 -17 581
rect 163 547 175 581
rect 355 547 367 581
rect 547 547 559 581
rect 739 547 751 581
rect 931 547 943 581
rect 1123 547 1135 581
rect -1181 541 -1123 547
rect -989 541 -931 547
rect -797 541 -739 547
rect -605 541 -547 547
rect -413 541 -355 547
rect -221 541 -163 547
rect -29 541 29 547
rect 163 541 221 547
rect 355 541 413 547
rect 547 541 605 547
rect 739 541 797 547
rect 931 541 989 547
rect 1123 541 1181 547
rect -1085 71 -1027 77
rect -893 71 -835 77
rect -701 71 -643 77
rect -509 71 -451 77
rect -317 71 -259 77
rect -125 71 -67 77
rect 67 71 125 77
rect 259 71 317 77
rect 451 71 509 77
rect 643 71 701 77
rect 835 71 893 77
rect 1027 71 1085 77
rect -1085 37 -1073 71
rect -893 37 -881 71
rect -701 37 -689 71
rect -509 37 -497 71
rect -317 37 -305 71
rect -125 37 -113 71
rect 67 37 79 71
rect 259 37 271 71
rect 451 37 463 71
rect 643 37 655 71
rect 835 37 847 71
rect 1027 37 1039 71
rect -1085 31 -1027 37
rect -893 31 -835 37
rect -701 31 -643 37
rect -509 31 -451 37
rect -317 31 -259 37
rect -125 31 -67 37
rect 67 31 125 37
rect 259 31 317 37
rect 451 31 509 37
rect 643 31 701 37
rect 835 31 893 37
rect 1027 31 1085 37
rect -1085 -37 -1027 -31
rect -893 -37 -835 -31
rect -701 -37 -643 -31
rect -509 -37 -451 -31
rect -317 -37 -259 -31
rect -125 -37 -67 -31
rect 67 -37 125 -31
rect 259 -37 317 -31
rect 451 -37 509 -31
rect 643 -37 701 -31
rect 835 -37 893 -31
rect 1027 -37 1085 -31
rect -1085 -71 -1073 -37
rect -893 -71 -881 -37
rect -701 -71 -689 -37
rect -509 -71 -497 -37
rect -317 -71 -305 -37
rect -125 -71 -113 -37
rect 67 -71 79 -37
rect 259 -71 271 -37
rect 451 -71 463 -37
rect 643 -71 655 -37
rect 835 -71 847 -37
rect 1027 -71 1039 -37
rect -1085 -77 -1027 -71
rect -893 -77 -835 -71
rect -701 -77 -643 -71
rect -509 -77 -451 -71
rect -317 -77 -259 -71
rect -125 -77 -67 -71
rect 67 -77 125 -71
rect 259 -77 317 -71
rect 451 -77 509 -71
rect 643 -77 701 -71
rect 835 -77 893 -71
rect 1027 -77 1085 -71
rect -1181 -547 -1123 -541
rect -989 -547 -931 -541
rect -797 -547 -739 -541
rect -605 -547 -547 -541
rect -413 -547 -355 -541
rect -221 -547 -163 -541
rect -29 -547 29 -541
rect 163 -547 221 -541
rect 355 -547 413 -541
rect 547 -547 605 -541
rect 739 -547 797 -541
rect 931 -547 989 -541
rect 1123 -547 1181 -541
rect -1181 -581 -1169 -547
rect -989 -581 -977 -547
rect -797 -581 -785 -547
rect -605 -581 -593 -547
rect -413 -581 -401 -547
rect -221 -581 -209 -547
rect -29 -581 -17 -547
rect 163 -581 175 -547
rect 355 -581 367 -547
rect 547 -581 559 -547
rect 739 -581 751 -547
rect 931 -581 943 -547
rect 1123 -581 1135 -547
rect -1181 -587 -1123 -581
rect -989 -587 -931 -581
rect -797 -587 -739 -581
rect -605 -587 -547 -581
rect -413 -587 -355 -581
rect -221 -587 -163 -581
rect -29 -587 29 -581
rect 163 -587 221 -581
rect 355 -587 413 -581
rect 547 -587 605 -581
rect 739 -587 797 -581
rect 931 -587 989 -581
rect 1123 -587 1181 -581
<< pwell >>
rect -1367 -719 1367 719
<< nmos >>
rect -1167 109 -1137 509
rect -1071 109 -1041 509
rect -975 109 -945 509
rect -879 109 -849 509
rect -783 109 -753 509
rect -687 109 -657 509
rect -591 109 -561 509
rect -495 109 -465 509
rect -399 109 -369 509
rect -303 109 -273 509
rect -207 109 -177 509
rect -111 109 -81 509
rect -15 109 15 509
rect 81 109 111 509
rect 177 109 207 509
rect 273 109 303 509
rect 369 109 399 509
rect 465 109 495 509
rect 561 109 591 509
rect 657 109 687 509
rect 753 109 783 509
rect 849 109 879 509
rect 945 109 975 509
rect 1041 109 1071 509
rect 1137 109 1167 509
rect -1167 -509 -1137 -109
rect -1071 -509 -1041 -109
rect -975 -509 -945 -109
rect -879 -509 -849 -109
rect -783 -509 -753 -109
rect -687 -509 -657 -109
rect -591 -509 -561 -109
rect -495 -509 -465 -109
rect -399 -509 -369 -109
rect -303 -509 -273 -109
rect -207 -509 -177 -109
rect -111 -509 -81 -109
rect -15 -509 15 -109
rect 81 -509 111 -109
rect 177 -509 207 -109
rect 273 -509 303 -109
rect 369 -509 399 -109
rect 465 -509 495 -109
rect 561 -509 591 -109
rect 657 -509 687 -109
rect 753 -509 783 -109
rect 849 -509 879 -109
rect 945 -509 975 -109
rect 1041 -509 1071 -109
rect 1137 -509 1167 -109
<< ndiff >>
rect -1229 497 -1167 509
rect -1229 121 -1217 497
rect -1183 121 -1167 497
rect -1229 109 -1167 121
rect -1137 497 -1071 509
rect -1137 121 -1121 497
rect -1087 121 -1071 497
rect -1137 109 -1071 121
rect -1041 497 -975 509
rect -1041 121 -1025 497
rect -991 121 -975 497
rect -1041 109 -975 121
rect -945 497 -879 509
rect -945 121 -929 497
rect -895 121 -879 497
rect -945 109 -879 121
rect -849 497 -783 509
rect -849 121 -833 497
rect -799 121 -783 497
rect -849 109 -783 121
rect -753 497 -687 509
rect -753 121 -737 497
rect -703 121 -687 497
rect -753 109 -687 121
rect -657 497 -591 509
rect -657 121 -641 497
rect -607 121 -591 497
rect -657 109 -591 121
rect -561 497 -495 509
rect -561 121 -545 497
rect -511 121 -495 497
rect -561 109 -495 121
rect -465 497 -399 509
rect -465 121 -449 497
rect -415 121 -399 497
rect -465 109 -399 121
rect -369 497 -303 509
rect -369 121 -353 497
rect -319 121 -303 497
rect -369 109 -303 121
rect -273 497 -207 509
rect -273 121 -257 497
rect -223 121 -207 497
rect -273 109 -207 121
rect -177 497 -111 509
rect -177 121 -161 497
rect -127 121 -111 497
rect -177 109 -111 121
rect -81 497 -15 509
rect -81 121 -65 497
rect -31 121 -15 497
rect -81 109 -15 121
rect 15 497 81 509
rect 15 121 31 497
rect 65 121 81 497
rect 15 109 81 121
rect 111 497 177 509
rect 111 121 127 497
rect 161 121 177 497
rect 111 109 177 121
rect 207 497 273 509
rect 207 121 223 497
rect 257 121 273 497
rect 207 109 273 121
rect 303 497 369 509
rect 303 121 319 497
rect 353 121 369 497
rect 303 109 369 121
rect 399 497 465 509
rect 399 121 415 497
rect 449 121 465 497
rect 399 109 465 121
rect 495 497 561 509
rect 495 121 511 497
rect 545 121 561 497
rect 495 109 561 121
rect 591 497 657 509
rect 591 121 607 497
rect 641 121 657 497
rect 591 109 657 121
rect 687 497 753 509
rect 687 121 703 497
rect 737 121 753 497
rect 687 109 753 121
rect 783 497 849 509
rect 783 121 799 497
rect 833 121 849 497
rect 783 109 849 121
rect 879 497 945 509
rect 879 121 895 497
rect 929 121 945 497
rect 879 109 945 121
rect 975 497 1041 509
rect 975 121 991 497
rect 1025 121 1041 497
rect 975 109 1041 121
rect 1071 497 1137 509
rect 1071 121 1087 497
rect 1121 121 1137 497
rect 1071 109 1137 121
rect 1167 497 1229 509
rect 1167 121 1183 497
rect 1217 121 1229 497
rect 1167 109 1229 121
rect -1229 -121 -1167 -109
rect -1229 -497 -1217 -121
rect -1183 -497 -1167 -121
rect -1229 -509 -1167 -497
rect -1137 -121 -1071 -109
rect -1137 -497 -1121 -121
rect -1087 -497 -1071 -121
rect -1137 -509 -1071 -497
rect -1041 -121 -975 -109
rect -1041 -497 -1025 -121
rect -991 -497 -975 -121
rect -1041 -509 -975 -497
rect -945 -121 -879 -109
rect -945 -497 -929 -121
rect -895 -497 -879 -121
rect -945 -509 -879 -497
rect -849 -121 -783 -109
rect -849 -497 -833 -121
rect -799 -497 -783 -121
rect -849 -509 -783 -497
rect -753 -121 -687 -109
rect -753 -497 -737 -121
rect -703 -497 -687 -121
rect -753 -509 -687 -497
rect -657 -121 -591 -109
rect -657 -497 -641 -121
rect -607 -497 -591 -121
rect -657 -509 -591 -497
rect -561 -121 -495 -109
rect -561 -497 -545 -121
rect -511 -497 -495 -121
rect -561 -509 -495 -497
rect -465 -121 -399 -109
rect -465 -497 -449 -121
rect -415 -497 -399 -121
rect -465 -509 -399 -497
rect -369 -121 -303 -109
rect -369 -497 -353 -121
rect -319 -497 -303 -121
rect -369 -509 -303 -497
rect -273 -121 -207 -109
rect -273 -497 -257 -121
rect -223 -497 -207 -121
rect -273 -509 -207 -497
rect -177 -121 -111 -109
rect -177 -497 -161 -121
rect -127 -497 -111 -121
rect -177 -509 -111 -497
rect -81 -121 -15 -109
rect -81 -497 -65 -121
rect -31 -497 -15 -121
rect -81 -509 -15 -497
rect 15 -121 81 -109
rect 15 -497 31 -121
rect 65 -497 81 -121
rect 15 -509 81 -497
rect 111 -121 177 -109
rect 111 -497 127 -121
rect 161 -497 177 -121
rect 111 -509 177 -497
rect 207 -121 273 -109
rect 207 -497 223 -121
rect 257 -497 273 -121
rect 207 -509 273 -497
rect 303 -121 369 -109
rect 303 -497 319 -121
rect 353 -497 369 -121
rect 303 -509 369 -497
rect 399 -121 465 -109
rect 399 -497 415 -121
rect 449 -497 465 -121
rect 399 -509 465 -497
rect 495 -121 561 -109
rect 495 -497 511 -121
rect 545 -497 561 -121
rect 495 -509 561 -497
rect 591 -121 657 -109
rect 591 -497 607 -121
rect 641 -497 657 -121
rect 591 -509 657 -497
rect 687 -121 753 -109
rect 687 -497 703 -121
rect 737 -497 753 -121
rect 687 -509 753 -497
rect 783 -121 849 -109
rect 783 -497 799 -121
rect 833 -497 849 -121
rect 783 -509 849 -497
rect 879 -121 945 -109
rect 879 -497 895 -121
rect 929 -497 945 -121
rect 879 -509 945 -497
rect 975 -121 1041 -109
rect 975 -497 991 -121
rect 1025 -497 1041 -121
rect 975 -509 1041 -497
rect 1071 -121 1137 -109
rect 1071 -497 1087 -121
rect 1121 -497 1137 -121
rect 1071 -509 1137 -497
rect 1167 -121 1229 -109
rect 1167 -497 1183 -121
rect 1217 -497 1229 -121
rect 1167 -509 1229 -497
<< ndiffc >>
rect -1217 121 -1183 497
rect -1121 121 -1087 497
rect -1025 121 -991 497
rect -929 121 -895 497
rect -833 121 -799 497
rect -737 121 -703 497
rect -641 121 -607 497
rect -545 121 -511 497
rect -449 121 -415 497
rect -353 121 -319 497
rect -257 121 -223 497
rect -161 121 -127 497
rect -65 121 -31 497
rect 31 121 65 497
rect 127 121 161 497
rect 223 121 257 497
rect 319 121 353 497
rect 415 121 449 497
rect 511 121 545 497
rect 607 121 641 497
rect 703 121 737 497
rect 799 121 833 497
rect 895 121 929 497
rect 991 121 1025 497
rect 1087 121 1121 497
rect 1183 121 1217 497
rect -1217 -497 -1183 -121
rect -1121 -497 -1087 -121
rect -1025 -497 -991 -121
rect -929 -497 -895 -121
rect -833 -497 -799 -121
rect -737 -497 -703 -121
rect -641 -497 -607 -121
rect -545 -497 -511 -121
rect -449 -497 -415 -121
rect -353 -497 -319 -121
rect -257 -497 -223 -121
rect -161 -497 -127 -121
rect -65 -497 -31 -121
rect 31 -497 65 -121
rect 127 -497 161 -121
rect 223 -497 257 -121
rect 319 -497 353 -121
rect 415 -497 449 -121
rect 511 -497 545 -121
rect 607 -497 641 -121
rect 703 -497 737 -121
rect 799 -497 833 -121
rect 895 -497 929 -121
rect 991 -497 1025 -121
rect 1087 -497 1121 -121
rect 1183 -497 1217 -121
<< psubdiff >>
rect -1331 649 -1235 683
rect 1235 649 1331 683
rect -1331 587 -1297 649
rect 1297 587 1331 649
rect -1331 -649 -1297 -587
rect 1297 -649 1331 -587
rect -1331 -683 -1235 -649
rect 1235 -683 1331 -649
<< psubdiffcont >>
rect -1235 649 1235 683
rect -1331 -587 -1297 587
rect 1297 -587 1331 587
rect -1235 -683 1235 -649
<< poly >>
rect -1185 581 -1119 597
rect -1185 547 -1169 581
rect -1135 547 -1119 581
rect -1185 531 -1119 547
rect -993 581 -927 597
rect -993 547 -977 581
rect -943 547 -927 581
rect -1167 509 -1137 531
rect -1071 509 -1041 535
rect -993 531 -927 547
rect -801 581 -735 597
rect -801 547 -785 581
rect -751 547 -735 581
rect -975 509 -945 531
rect -879 509 -849 535
rect -801 531 -735 547
rect -609 581 -543 597
rect -609 547 -593 581
rect -559 547 -543 581
rect -783 509 -753 531
rect -687 509 -657 535
rect -609 531 -543 547
rect -417 581 -351 597
rect -417 547 -401 581
rect -367 547 -351 581
rect -591 509 -561 531
rect -495 509 -465 535
rect -417 531 -351 547
rect -225 581 -159 597
rect -225 547 -209 581
rect -175 547 -159 581
rect -399 509 -369 531
rect -303 509 -273 535
rect -225 531 -159 547
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -207 509 -177 531
rect -111 509 -81 535
rect -33 531 33 547
rect 159 581 225 597
rect 159 547 175 581
rect 209 547 225 581
rect -15 509 15 531
rect 81 509 111 535
rect 159 531 225 547
rect 351 581 417 597
rect 351 547 367 581
rect 401 547 417 581
rect 177 509 207 531
rect 273 509 303 535
rect 351 531 417 547
rect 543 581 609 597
rect 543 547 559 581
rect 593 547 609 581
rect 369 509 399 531
rect 465 509 495 535
rect 543 531 609 547
rect 735 581 801 597
rect 735 547 751 581
rect 785 547 801 581
rect 561 509 591 531
rect 657 509 687 535
rect 735 531 801 547
rect 927 581 993 597
rect 927 547 943 581
rect 977 547 993 581
rect 753 509 783 531
rect 849 509 879 535
rect 927 531 993 547
rect 1119 581 1185 597
rect 1119 547 1135 581
rect 1169 547 1185 581
rect 945 509 975 531
rect 1041 509 1071 535
rect 1119 531 1185 547
rect 1137 509 1167 531
rect -1167 83 -1137 109
rect -1071 87 -1041 109
rect -1089 71 -1023 87
rect -975 83 -945 109
rect -879 87 -849 109
rect -1089 37 -1073 71
rect -1039 37 -1023 71
rect -1089 21 -1023 37
rect -897 71 -831 87
rect -783 83 -753 109
rect -687 87 -657 109
rect -897 37 -881 71
rect -847 37 -831 71
rect -897 21 -831 37
rect -705 71 -639 87
rect -591 83 -561 109
rect -495 87 -465 109
rect -705 37 -689 71
rect -655 37 -639 71
rect -705 21 -639 37
rect -513 71 -447 87
rect -399 83 -369 109
rect -303 87 -273 109
rect -513 37 -497 71
rect -463 37 -447 71
rect -513 21 -447 37
rect -321 71 -255 87
rect -207 83 -177 109
rect -111 87 -81 109
rect -321 37 -305 71
rect -271 37 -255 71
rect -321 21 -255 37
rect -129 71 -63 87
rect -15 83 15 109
rect 81 87 111 109
rect -129 37 -113 71
rect -79 37 -63 71
rect -129 21 -63 37
rect 63 71 129 87
rect 177 83 207 109
rect 273 87 303 109
rect 63 37 79 71
rect 113 37 129 71
rect 63 21 129 37
rect 255 71 321 87
rect 369 83 399 109
rect 465 87 495 109
rect 255 37 271 71
rect 305 37 321 71
rect 255 21 321 37
rect 447 71 513 87
rect 561 83 591 109
rect 657 87 687 109
rect 447 37 463 71
rect 497 37 513 71
rect 447 21 513 37
rect 639 71 705 87
rect 753 83 783 109
rect 849 87 879 109
rect 639 37 655 71
rect 689 37 705 71
rect 639 21 705 37
rect 831 71 897 87
rect 945 83 975 109
rect 1041 87 1071 109
rect 831 37 847 71
rect 881 37 897 71
rect 831 21 897 37
rect 1023 71 1089 87
rect 1137 83 1167 109
rect 1023 37 1039 71
rect 1073 37 1089 71
rect 1023 21 1089 37
rect -1089 -37 -1023 -21
rect -1089 -71 -1073 -37
rect -1039 -71 -1023 -37
rect -1167 -109 -1137 -83
rect -1089 -87 -1023 -71
rect -897 -37 -831 -21
rect -897 -71 -881 -37
rect -847 -71 -831 -37
rect -1071 -109 -1041 -87
rect -975 -109 -945 -83
rect -897 -87 -831 -71
rect -705 -37 -639 -21
rect -705 -71 -689 -37
rect -655 -71 -639 -37
rect -879 -109 -849 -87
rect -783 -109 -753 -83
rect -705 -87 -639 -71
rect -513 -37 -447 -21
rect -513 -71 -497 -37
rect -463 -71 -447 -37
rect -687 -109 -657 -87
rect -591 -109 -561 -83
rect -513 -87 -447 -71
rect -321 -37 -255 -21
rect -321 -71 -305 -37
rect -271 -71 -255 -37
rect -495 -109 -465 -87
rect -399 -109 -369 -83
rect -321 -87 -255 -71
rect -129 -37 -63 -21
rect -129 -71 -113 -37
rect -79 -71 -63 -37
rect -303 -109 -273 -87
rect -207 -109 -177 -83
rect -129 -87 -63 -71
rect 63 -37 129 -21
rect 63 -71 79 -37
rect 113 -71 129 -37
rect -111 -109 -81 -87
rect -15 -109 15 -83
rect 63 -87 129 -71
rect 255 -37 321 -21
rect 255 -71 271 -37
rect 305 -71 321 -37
rect 81 -109 111 -87
rect 177 -109 207 -83
rect 255 -87 321 -71
rect 447 -37 513 -21
rect 447 -71 463 -37
rect 497 -71 513 -37
rect 273 -109 303 -87
rect 369 -109 399 -83
rect 447 -87 513 -71
rect 639 -37 705 -21
rect 639 -71 655 -37
rect 689 -71 705 -37
rect 465 -109 495 -87
rect 561 -109 591 -83
rect 639 -87 705 -71
rect 831 -37 897 -21
rect 831 -71 847 -37
rect 881 -71 897 -37
rect 657 -109 687 -87
rect 753 -109 783 -83
rect 831 -87 897 -71
rect 1023 -37 1089 -21
rect 1023 -71 1039 -37
rect 1073 -71 1089 -37
rect 849 -109 879 -87
rect 945 -109 975 -83
rect 1023 -87 1089 -71
rect 1041 -109 1071 -87
rect 1137 -109 1167 -83
rect -1167 -531 -1137 -509
rect -1185 -547 -1119 -531
rect -1071 -535 -1041 -509
rect -975 -531 -945 -509
rect -1185 -581 -1169 -547
rect -1135 -581 -1119 -547
rect -1185 -597 -1119 -581
rect -993 -547 -927 -531
rect -879 -535 -849 -509
rect -783 -531 -753 -509
rect -993 -581 -977 -547
rect -943 -581 -927 -547
rect -993 -597 -927 -581
rect -801 -547 -735 -531
rect -687 -535 -657 -509
rect -591 -531 -561 -509
rect -801 -581 -785 -547
rect -751 -581 -735 -547
rect -801 -597 -735 -581
rect -609 -547 -543 -531
rect -495 -535 -465 -509
rect -399 -531 -369 -509
rect -609 -581 -593 -547
rect -559 -581 -543 -547
rect -609 -597 -543 -581
rect -417 -547 -351 -531
rect -303 -535 -273 -509
rect -207 -531 -177 -509
rect -417 -581 -401 -547
rect -367 -581 -351 -547
rect -417 -597 -351 -581
rect -225 -547 -159 -531
rect -111 -535 -81 -509
rect -15 -531 15 -509
rect -225 -581 -209 -547
rect -175 -581 -159 -547
rect -225 -597 -159 -581
rect -33 -547 33 -531
rect 81 -535 111 -509
rect 177 -531 207 -509
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
rect 159 -547 225 -531
rect 273 -535 303 -509
rect 369 -531 399 -509
rect 159 -581 175 -547
rect 209 -581 225 -547
rect 159 -597 225 -581
rect 351 -547 417 -531
rect 465 -535 495 -509
rect 561 -531 591 -509
rect 351 -581 367 -547
rect 401 -581 417 -547
rect 351 -597 417 -581
rect 543 -547 609 -531
rect 657 -535 687 -509
rect 753 -531 783 -509
rect 543 -581 559 -547
rect 593 -581 609 -547
rect 543 -597 609 -581
rect 735 -547 801 -531
rect 849 -535 879 -509
rect 945 -531 975 -509
rect 735 -581 751 -547
rect 785 -581 801 -547
rect 735 -597 801 -581
rect 927 -547 993 -531
rect 1041 -535 1071 -509
rect 1137 -531 1167 -509
rect 927 -581 943 -547
rect 977 -581 993 -547
rect 927 -597 993 -581
rect 1119 -547 1185 -531
rect 1119 -581 1135 -547
rect 1169 -581 1185 -547
rect 1119 -597 1185 -581
<< polycont >>
rect -1169 547 -1135 581
rect -977 547 -943 581
rect -785 547 -751 581
rect -593 547 -559 581
rect -401 547 -367 581
rect -209 547 -175 581
rect -17 547 17 581
rect 175 547 209 581
rect 367 547 401 581
rect 559 547 593 581
rect 751 547 785 581
rect 943 547 977 581
rect 1135 547 1169 581
rect -1073 37 -1039 71
rect -881 37 -847 71
rect -689 37 -655 71
rect -497 37 -463 71
rect -305 37 -271 71
rect -113 37 -79 71
rect 79 37 113 71
rect 271 37 305 71
rect 463 37 497 71
rect 655 37 689 71
rect 847 37 881 71
rect 1039 37 1073 71
rect -1073 -71 -1039 -37
rect -881 -71 -847 -37
rect -689 -71 -655 -37
rect -497 -71 -463 -37
rect -305 -71 -271 -37
rect -113 -71 -79 -37
rect 79 -71 113 -37
rect 271 -71 305 -37
rect 463 -71 497 -37
rect 655 -71 689 -37
rect 847 -71 881 -37
rect 1039 -71 1073 -37
rect -1169 -581 -1135 -547
rect -977 -581 -943 -547
rect -785 -581 -751 -547
rect -593 -581 -559 -547
rect -401 -581 -367 -547
rect -209 -581 -175 -547
rect -17 -581 17 -547
rect 175 -581 209 -547
rect 367 -581 401 -547
rect 559 -581 593 -547
rect 751 -581 785 -547
rect 943 -581 977 -547
rect 1135 -581 1169 -547
<< locali >>
rect -1331 649 -1235 683
rect 1235 649 1331 683
rect -1331 587 -1297 649
rect 1297 587 1331 649
rect -1185 547 -1169 581
rect -1135 547 -1119 581
rect -993 547 -977 581
rect -943 547 -927 581
rect -801 547 -785 581
rect -751 547 -735 581
rect -609 547 -593 581
rect -559 547 -543 581
rect -417 547 -401 581
rect -367 547 -351 581
rect -225 547 -209 581
rect -175 547 -159 581
rect -33 547 -17 581
rect 17 547 33 581
rect 159 547 175 581
rect 209 547 225 581
rect 351 547 367 581
rect 401 547 417 581
rect 543 547 559 581
rect 593 547 609 581
rect 735 547 751 581
rect 785 547 801 581
rect 927 547 943 581
rect 977 547 993 581
rect 1119 547 1135 581
rect 1169 547 1185 581
rect -1217 497 -1183 513
rect -1217 105 -1183 121
rect -1121 497 -1087 513
rect -1121 105 -1087 121
rect -1025 497 -991 513
rect -1025 105 -991 121
rect -929 497 -895 513
rect -929 105 -895 121
rect -833 497 -799 513
rect -833 105 -799 121
rect -737 497 -703 513
rect -737 105 -703 121
rect -641 497 -607 513
rect -641 105 -607 121
rect -545 497 -511 513
rect -545 105 -511 121
rect -449 497 -415 513
rect -449 105 -415 121
rect -353 497 -319 513
rect -353 105 -319 121
rect -257 497 -223 513
rect -257 105 -223 121
rect -161 497 -127 513
rect -161 105 -127 121
rect -65 497 -31 513
rect -65 105 -31 121
rect 31 497 65 513
rect 31 105 65 121
rect 127 497 161 513
rect 127 105 161 121
rect 223 497 257 513
rect 223 105 257 121
rect 319 497 353 513
rect 319 105 353 121
rect 415 497 449 513
rect 415 105 449 121
rect 511 497 545 513
rect 511 105 545 121
rect 607 497 641 513
rect 607 105 641 121
rect 703 497 737 513
rect 703 105 737 121
rect 799 497 833 513
rect 799 105 833 121
rect 895 497 929 513
rect 895 105 929 121
rect 991 497 1025 513
rect 991 105 1025 121
rect 1087 497 1121 513
rect 1087 105 1121 121
rect 1183 497 1217 513
rect 1183 105 1217 121
rect -1089 37 -1073 71
rect -1039 37 -1023 71
rect -897 37 -881 71
rect -847 37 -831 71
rect -705 37 -689 71
rect -655 37 -639 71
rect -513 37 -497 71
rect -463 37 -447 71
rect -321 37 -305 71
rect -271 37 -255 71
rect -129 37 -113 71
rect -79 37 -63 71
rect 63 37 79 71
rect 113 37 129 71
rect 255 37 271 71
rect 305 37 321 71
rect 447 37 463 71
rect 497 37 513 71
rect 639 37 655 71
rect 689 37 705 71
rect 831 37 847 71
rect 881 37 897 71
rect 1023 37 1039 71
rect 1073 37 1089 71
rect -1089 -71 -1073 -37
rect -1039 -71 -1023 -37
rect -897 -71 -881 -37
rect -847 -71 -831 -37
rect -705 -71 -689 -37
rect -655 -71 -639 -37
rect -513 -71 -497 -37
rect -463 -71 -447 -37
rect -321 -71 -305 -37
rect -271 -71 -255 -37
rect -129 -71 -113 -37
rect -79 -71 -63 -37
rect 63 -71 79 -37
rect 113 -71 129 -37
rect 255 -71 271 -37
rect 305 -71 321 -37
rect 447 -71 463 -37
rect 497 -71 513 -37
rect 639 -71 655 -37
rect 689 -71 705 -37
rect 831 -71 847 -37
rect 881 -71 897 -37
rect 1023 -71 1039 -37
rect 1073 -71 1089 -37
rect -1217 -121 -1183 -105
rect -1217 -513 -1183 -497
rect -1121 -121 -1087 -105
rect -1121 -513 -1087 -497
rect -1025 -121 -991 -105
rect -1025 -513 -991 -497
rect -929 -121 -895 -105
rect -929 -513 -895 -497
rect -833 -121 -799 -105
rect -833 -513 -799 -497
rect -737 -121 -703 -105
rect -737 -513 -703 -497
rect -641 -121 -607 -105
rect -641 -513 -607 -497
rect -545 -121 -511 -105
rect -545 -513 -511 -497
rect -449 -121 -415 -105
rect -449 -513 -415 -497
rect -353 -121 -319 -105
rect -353 -513 -319 -497
rect -257 -121 -223 -105
rect -257 -513 -223 -497
rect -161 -121 -127 -105
rect -161 -513 -127 -497
rect -65 -121 -31 -105
rect -65 -513 -31 -497
rect 31 -121 65 -105
rect 31 -513 65 -497
rect 127 -121 161 -105
rect 127 -513 161 -497
rect 223 -121 257 -105
rect 223 -513 257 -497
rect 319 -121 353 -105
rect 319 -513 353 -497
rect 415 -121 449 -105
rect 415 -513 449 -497
rect 511 -121 545 -105
rect 511 -513 545 -497
rect 607 -121 641 -105
rect 607 -513 641 -497
rect 703 -121 737 -105
rect 703 -513 737 -497
rect 799 -121 833 -105
rect 799 -513 833 -497
rect 895 -121 929 -105
rect 895 -513 929 -497
rect 991 -121 1025 -105
rect 991 -513 1025 -497
rect 1087 -121 1121 -105
rect 1087 -513 1121 -497
rect 1183 -121 1217 -105
rect 1183 -513 1217 -497
rect -1185 -581 -1169 -547
rect -1135 -581 -1119 -547
rect -993 -581 -977 -547
rect -943 -581 -927 -547
rect -801 -581 -785 -547
rect -751 -581 -735 -547
rect -609 -581 -593 -547
rect -559 -581 -543 -547
rect -417 -581 -401 -547
rect -367 -581 -351 -547
rect -225 -581 -209 -547
rect -175 -581 -159 -547
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect 159 -581 175 -547
rect 209 -581 225 -547
rect 351 -581 367 -547
rect 401 -581 417 -547
rect 543 -581 559 -547
rect 593 -581 609 -547
rect 735 -581 751 -547
rect 785 -581 801 -547
rect 927 -581 943 -547
rect 977 -581 993 -547
rect 1119 -581 1135 -547
rect 1169 -581 1185 -547
rect -1331 -649 -1297 -587
rect 1297 -649 1331 -587
rect -1331 -683 -1235 -649
rect 1235 -683 1331 -649
<< viali >>
rect -1169 547 -1135 581
rect -977 547 -943 581
rect -785 547 -751 581
rect -593 547 -559 581
rect -401 547 -367 581
rect -209 547 -175 581
rect -17 547 17 581
rect 175 547 209 581
rect 367 547 401 581
rect 559 547 593 581
rect 751 547 785 581
rect 943 547 977 581
rect 1135 547 1169 581
rect -1217 121 -1183 497
rect -1121 121 -1087 497
rect -1025 121 -991 497
rect -929 121 -895 497
rect -833 121 -799 497
rect -737 121 -703 497
rect -641 121 -607 497
rect -545 121 -511 497
rect -449 121 -415 497
rect -353 121 -319 497
rect -257 121 -223 497
rect -161 121 -127 497
rect -65 121 -31 497
rect 31 121 65 497
rect 127 121 161 497
rect 223 121 257 497
rect 319 121 353 497
rect 415 121 449 497
rect 511 121 545 497
rect 607 121 641 497
rect 703 121 737 497
rect 799 121 833 497
rect 895 121 929 497
rect 991 121 1025 497
rect 1087 121 1121 497
rect 1183 121 1217 497
rect -1073 37 -1039 71
rect -881 37 -847 71
rect -689 37 -655 71
rect -497 37 -463 71
rect -305 37 -271 71
rect -113 37 -79 71
rect 79 37 113 71
rect 271 37 305 71
rect 463 37 497 71
rect 655 37 689 71
rect 847 37 881 71
rect 1039 37 1073 71
rect -1073 -71 -1039 -37
rect -881 -71 -847 -37
rect -689 -71 -655 -37
rect -497 -71 -463 -37
rect -305 -71 -271 -37
rect -113 -71 -79 -37
rect 79 -71 113 -37
rect 271 -71 305 -37
rect 463 -71 497 -37
rect 655 -71 689 -37
rect 847 -71 881 -37
rect 1039 -71 1073 -37
rect -1217 -497 -1183 -121
rect -1121 -497 -1087 -121
rect -1025 -497 -991 -121
rect -929 -497 -895 -121
rect -833 -497 -799 -121
rect -737 -497 -703 -121
rect -641 -497 -607 -121
rect -545 -497 -511 -121
rect -449 -497 -415 -121
rect -353 -497 -319 -121
rect -257 -497 -223 -121
rect -161 -497 -127 -121
rect -65 -497 -31 -121
rect 31 -497 65 -121
rect 127 -497 161 -121
rect 223 -497 257 -121
rect 319 -497 353 -121
rect 415 -497 449 -121
rect 511 -497 545 -121
rect 607 -497 641 -121
rect 703 -497 737 -121
rect 799 -497 833 -121
rect 895 -497 929 -121
rect 991 -497 1025 -121
rect 1087 -497 1121 -121
rect 1183 -497 1217 -121
rect -1169 -581 -1135 -547
rect -977 -581 -943 -547
rect -785 -581 -751 -547
rect -593 -581 -559 -547
rect -401 -581 -367 -547
rect -209 -581 -175 -547
rect -17 -581 17 -547
rect 175 -581 209 -547
rect 367 -581 401 -547
rect 559 -581 593 -547
rect 751 -581 785 -547
rect 943 -581 977 -547
rect 1135 -581 1169 -547
<< metal1 >>
rect -1181 581 -1123 587
rect -1181 547 -1169 581
rect -1135 547 -1123 581
rect -1181 541 -1123 547
rect -989 581 -931 587
rect -989 547 -977 581
rect -943 547 -931 581
rect -989 541 -931 547
rect -797 581 -739 587
rect -797 547 -785 581
rect -751 547 -739 581
rect -797 541 -739 547
rect -605 581 -547 587
rect -605 547 -593 581
rect -559 547 -547 581
rect -605 541 -547 547
rect -413 581 -355 587
rect -413 547 -401 581
rect -367 547 -355 581
rect -413 541 -355 547
rect -221 581 -163 587
rect -221 547 -209 581
rect -175 547 -163 581
rect -221 541 -163 547
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect 163 581 221 587
rect 163 547 175 581
rect 209 547 221 581
rect 163 541 221 547
rect 355 581 413 587
rect 355 547 367 581
rect 401 547 413 581
rect 355 541 413 547
rect 547 581 605 587
rect 547 547 559 581
rect 593 547 605 581
rect 547 541 605 547
rect 739 581 797 587
rect 739 547 751 581
rect 785 547 797 581
rect 739 541 797 547
rect 931 581 989 587
rect 931 547 943 581
rect 977 547 989 581
rect 931 541 989 547
rect 1123 581 1181 587
rect 1123 547 1135 581
rect 1169 547 1181 581
rect 1123 541 1181 547
rect -1223 497 -1177 509
rect -1223 121 -1217 497
rect -1183 121 -1177 497
rect -1223 109 -1177 121
rect -1127 497 -1081 509
rect -1127 121 -1121 497
rect -1087 121 -1081 497
rect -1127 109 -1081 121
rect -1031 497 -985 509
rect -1031 121 -1025 497
rect -991 121 -985 497
rect -1031 109 -985 121
rect -935 497 -889 509
rect -935 121 -929 497
rect -895 121 -889 497
rect -935 109 -889 121
rect -839 497 -793 509
rect -839 121 -833 497
rect -799 121 -793 497
rect -839 109 -793 121
rect -743 497 -697 509
rect -743 121 -737 497
rect -703 121 -697 497
rect -743 109 -697 121
rect -647 497 -601 509
rect -647 121 -641 497
rect -607 121 -601 497
rect -647 109 -601 121
rect -551 497 -505 509
rect -551 121 -545 497
rect -511 121 -505 497
rect -551 109 -505 121
rect -455 497 -409 509
rect -455 121 -449 497
rect -415 121 -409 497
rect -455 109 -409 121
rect -359 497 -313 509
rect -359 121 -353 497
rect -319 121 -313 497
rect -359 109 -313 121
rect -263 497 -217 509
rect -263 121 -257 497
rect -223 121 -217 497
rect -263 109 -217 121
rect -167 497 -121 509
rect -167 121 -161 497
rect -127 121 -121 497
rect -167 109 -121 121
rect -71 497 -25 509
rect -71 121 -65 497
rect -31 121 -25 497
rect -71 109 -25 121
rect 25 497 71 509
rect 25 121 31 497
rect 65 121 71 497
rect 25 109 71 121
rect 121 497 167 509
rect 121 121 127 497
rect 161 121 167 497
rect 121 109 167 121
rect 217 497 263 509
rect 217 121 223 497
rect 257 121 263 497
rect 217 109 263 121
rect 313 497 359 509
rect 313 121 319 497
rect 353 121 359 497
rect 313 109 359 121
rect 409 497 455 509
rect 409 121 415 497
rect 449 121 455 497
rect 409 109 455 121
rect 505 497 551 509
rect 505 121 511 497
rect 545 121 551 497
rect 505 109 551 121
rect 601 497 647 509
rect 601 121 607 497
rect 641 121 647 497
rect 601 109 647 121
rect 697 497 743 509
rect 697 121 703 497
rect 737 121 743 497
rect 697 109 743 121
rect 793 497 839 509
rect 793 121 799 497
rect 833 121 839 497
rect 793 109 839 121
rect 889 497 935 509
rect 889 121 895 497
rect 929 121 935 497
rect 889 109 935 121
rect 985 497 1031 509
rect 985 121 991 497
rect 1025 121 1031 497
rect 985 109 1031 121
rect 1081 497 1127 509
rect 1081 121 1087 497
rect 1121 121 1127 497
rect 1081 109 1127 121
rect 1177 497 1223 509
rect 1177 121 1183 497
rect 1217 121 1223 497
rect 1177 109 1223 121
rect -1085 71 -1027 77
rect -1085 37 -1073 71
rect -1039 37 -1027 71
rect -1085 31 -1027 37
rect -893 71 -835 77
rect -893 37 -881 71
rect -847 37 -835 71
rect -893 31 -835 37
rect -701 71 -643 77
rect -701 37 -689 71
rect -655 37 -643 71
rect -701 31 -643 37
rect -509 71 -451 77
rect -509 37 -497 71
rect -463 37 -451 71
rect -509 31 -451 37
rect -317 71 -259 77
rect -317 37 -305 71
rect -271 37 -259 71
rect -317 31 -259 37
rect -125 71 -67 77
rect -125 37 -113 71
rect -79 37 -67 71
rect -125 31 -67 37
rect 67 71 125 77
rect 67 37 79 71
rect 113 37 125 71
rect 67 31 125 37
rect 259 71 317 77
rect 259 37 271 71
rect 305 37 317 71
rect 259 31 317 37
rect 451 71 509 77
rect 451 37 463 71
rect 497 37 509 71
rect 451 31 509 37
rect 643 71 701 77
rect 643 37 655 71
rect 689 37 701 71
rect 643 31 701 37
rect 835 71 893 77
rect 835 37 847 71
rect 881 37 893 71
rect 835 31 893 37
rect 1027 71 1085 77
rect 1027 37 1039 71
rect 1073 37 1085 71
rect 1027 31 1085 37
rect -1085 -37 -1027 -31
rect -1085 -71 -1073 -37
rect -1039 -71 -1027 -37
rect -1085 -77 -1027 -71
rect -893 -37 -835 -31
rect -893 -71 -881 -37
rect -847 -71 -835 -37
rect -893 -77 -835 -71
rect -701 -37 -643 -31
rect -701 -71 -689 -37
rect -655 -71 -643 -37
rect -701 -77 -643 -71
rect -509 -37 -451 -31
rect -509 -71 -497 -37
rect -463 -71 -451 -37
rect -509 -77 -451 -71
rect -317 -37 -259 -31
rect -317 -71 -305 -37
rect -271 -71 -259 -37
rect -317 -77 -259 -71
rect -125 -37 -67 -31
rect -125 -71 -113 -37
rect -79 -71 -67 -37
rect -125 -77 -67 -71
rect 67 -37 125 -31
rect 67 -71 79 -37
rect 113 -71 125 -37
rect 67 -77 125 -71
rect 259 -37 317 -31
rect 259 -71 271 -37
rect 305 -71 317 -37
rect 259 -77 317 -71
rect 451 -37 509 -31
rect 451 -71 463 -37
rect 497 -71 509 -37
rect 451 -77 509 -71
rect 643 -37 701 -31
rect 643 -71 655 -37
rect 689 -71 701 -37
rect 643 -77 701 -71
rect 835 -37 893 -31
rect 835 -71 847 -37
rect 881 -71 893 -37
rect 835 -77 893 -71
rect 1027 -37 1085 -31
rect 1027 -71 1039 -37
rect 1073 -71 1085 -37
rect 1027 -77 1085 -71
rect -1223 -121 -1177 -109
rect -1223 -497 -1217 -121
rect -1183 -497 -1177 -121
rect -1223 -509 -1177 -497
rect -1127 -121 -1081 -109
rect -1127 -497 -1121 -121
rect -1087 -497 -1081 -121
rect -1127 -509 -1081 -497
rect -1031 -121 -985 -109
rect -1031 -497 -1025 -121
rect -991 -497 -985 -121
rect -1031 -509 -985 -497
rect -935 -121 -889 -109
rect -935 -497 -929 -121
rect -895 -497 -889 -121
rect -935 -509 -889 -497
rect -839 -121 -793 -109
rect -839 -497 -833 -121
rect -799 -497 -793 -121
rect -839 -509 -793 -497
rect -743 -121 -697 -109
rect -743 -497 -737 -121
rect -703 -497 -697 -121
rect -743 -509 -697 -497
rect -647 -121 -601 -109
rect -647 -497 -641 -121
rect -607 -497 -601 -121
rect -647 -509 -601 -497
rect -551 -121 -505 -109
rect -551 -497 -545 -121
rect -511 -497 -505 -121
rect -551 -509 -505 -497
rect -455 -121 -409 -109
rect -455 -497 -449 -121
rect -415 -497 -409 -121
rect -455 -509 -409 -497
rect -359 -121 -313 -109
rect -359 -497 -353 -121
rect -319 -497 -313 -121
rect -359 -509 -313 -497
rect -263 -121 -217 -109
rect -263 -497 -257 -121
rect -223 -497 -217 -121
rect -263 -509 -217 -497
rect -167 -121 -121 -109
rect -167 -497 -161 -121
rect -127 -497 -121 -121
rect -167 -509 -121 -497
rect -71 -121 -25 -109
rect -71 -497 -65 -121
rect -31 -497 -25 -121
rect -71 -509 -25 -497
rect 25 -121 71 -109
rect 25 -497 31 -121
rect 65 -497 71 -121
rect 25 -509 71 -497
rect 121 -121 167 -109
rect 121 -497 127 -121
rect 161 -497 167 -121
rect 121 -509 167 -497
rect 217 -121 263 -109
rect 217 -497 223 -121
rect 257 -497 263 -121
rect 217 -509 263 -497
rect 313 -121 359 -109
rect 313 -497 319 -121
rect 353 -497 359 -121
rect 313 -509 359 -497
rect 409 -121 455 -109
rect 409 -497 415 -121
rect 449 -497 455 -121
rect 409 -509 455 -497
rect 505 -121 551 -109
rect 505 -497 511 -121
rect 545 -497 551 -121
rect 505 -509 551 -497
rect 601 -121 647 -109
rect 601 -497 607 -121
rect 641 -497 647 -121
rect 601 -509 647 -497
rect 697 -121 743 -109
rect 697 -497 703 -121
rect 737 -497 743 -121
rect 697 -509 743 -497
rect 793 -121 839 -109
rect 793 -497 799 -121
rect 833 -497 839 -121
rect 793 -509 839 -497
rect 889 -121 935 -109
rect 889 -497 895 -121
rect 929 -497 935 -121
rect 889 -509 935 -497
rect 985 -121 1031 -109
rect 985 -497 991 -121
rect 1025 -497 1031 -121
rect 985 -509 1031 -497
rect 1081 -121 1127 -109
rect 1081 -497 1087 -121
rect 1121 -497 1127 -121
rect 1081 -509 1127 -497
rect 1177 -121 1223 -109
rect 1177 -497 1183 -121
rect 1217 -497 1223 -121
rect 1177 -509 1223 -497
rect -1181 -547 -1123 -541
rect -1181 -581 -1169 -547
rect -1135 -581 -1123 -547
rect -1181 -587 -1123 -581
rect -989 -547 -931 -541
rect -989 -581 -977 -547
rect -943 -581 -931 -547
rect -989 -587 -931 -581
rect -797 -547 -739 -541
rect -797 -581 -785 -547
rect -751 -581 -739 -547
rect -797 -587 -739 -581
rect -605 -547 -547 -541
rect -605 -581 -593 -547
rect -559 -581 -547 -547
rect -605 -587 -547 -581
rect -413 -547 -355 -541
rect -413 -581 -401 -547
rect -367 -581 -355 -547
rect -413 -587 -355 -581
rect -221 -547 -163 -541
rect -221 -581 -209 -547
rect -175 -581 -163 -547
rect -221 -587 -163 -581
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
rect 163 -547 221 -541
rect 163 -581 175 -547
rect 209 -581 221 -547
rect 163 -587 221 -581
rect 355 -547 413 -541
rect 355 -581 367 -547
rect 401 -581 413 -547
rect 355 -587 413 -581
rect 547 -547 605 -541
rect 547 -581 559 -547
rect 593 -581 605 -547
rect 547 -587 605 -581
rect 739 -547 797 -541
rect 739 -581 751 -547
rect 785 -581 797 -547
rect 739 -587 797 -581
rect 931 -547 989 -541
rect 931 -581 943 -547
rect 977 -581 989 -547
rect 931 -587 989 -581
rect 1123 -547 1181 -541
rect 1123 -581 1135 -547
rect 1169 -581 1181 -547
rect 1123 -587 1181 -581
<< properties >>
string FIXED_BBOX -1314 -666 1314 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 2 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
