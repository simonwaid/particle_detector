magic
tech sky130A
magscale 1 2
timestamp 1646234887
<< pwell >>
rect -1431 -410 1431 410
<< nmos >>
rect -1235 -200 -1135 200
rect -1077 -200 -977 200
rect -919 -200 -819 200
rect -761 -200 -661 200
rect -603 -200 -503 200
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
rect 503 -200 603 200
rect 661 -200 761 200
rect 819 -200 919 200
rect 977 -200 1077 200
rect 1135 -200 1235 200
<< ndiff >>
rect -1293 188 -1235 200
rect -1293 -188 -1281 188
rect -1247 -188 -1235 188
rect -1293 -200 -1235 -188
rect -1135 188 -1077 200
rect -1135 -188 -1123 188
rect -1089 -188 -1077 188
rect -1135 -200 -1077 -188
rect -977 188 -919 200
rect -977 -188 -965 188
rect -931 -188 -919 188
rect -977 -200 -919 -188
rect -819 188 -761 200
rect -819 -188 -807 188
rect -773 -188 -761 188
rect -819 -200 -761 -188
rect -661 188 -603 200
rect -661 -188 -649 188
rect -615 -188 -603 188
rect -661 -200 -603 -188
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
rect 603 188 661 200
rect 603 -188 615 188
rect 649 -188 661 188
rect 603 -200 661 -188
rect 761 188 819 200
rect 761 -188 773 188
rect 807 -188 819 188
rect 761 -200 819 -188
rect 919 188 977 200
rect 919 -188 931 188
rect 965 -188 977 188
rect 919 -200 977 -188
rect 1077 188 1135 200
rect 1077 -188 1089 188
rect 1123 -188 1135 188
rect 1077 -200 1135 -188
rect 1235 188 1293 200
rect 1235 -188 1247 188
rect 1281 -188 1293 188
rect 1235 -200 1293 -188
<< ndiffc >>
rect -1281 -188 -1247 188
rect -1123 -188 -1089 188
rect -965 -188 -931 188
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect 931 -188 965 188
rect 1089 -188 1123 188
rect 1247 -188 1281 188
<< psubdiff >>
rect -1395 340 -1299 374
rect 1299 340 1395 374
rect -1395 278 -1361 340
rect 1361 278 1395 340
rect -1395 -340 -1361 -278
rect 1361 -340 1395 -278
rect -1395 -374 -1299 -340
rect 1299 -374 1395 -340
<< psubdiffcont >>
rect -1299 340 1299 374
rect -1395 -278 -1361 278
rect 1361 -278 1395 278
rect -1299 -374 1299 -340
<< poly >>
rect -1235 272 -1135 288
rect -1235 238 -1219 272
rect -1151 238 -1135 272
rect -1235 200 -1135 238
rect -1077 272 -977 288
rect -1077 238 -1061 272
rect -993 238 -977 272
rect -1077 200 -977 238
rect -919 272 -819 288
rect -919 238 -903 272
rect -835 238 -819 272
rect -919 200 -819 238
rect -761 272 -661 288
rect -761 238 -745 272
rect -677 238 -661 272
rect -761 200 -661 238
rect -603 272 -503 288
rect -603 238 -587 272
rect -519 238 -503 272
rect -603 200 -503 238
rect -445 272 -345 288
rect -445 238 -429 272
rect -361 238 -345 272
rect -445 200 -345 238
rect -287 272 -187 288
rect -287 238 -271 272
rect -203 238 -187 272
rect -287 200 -187 238
rect -129 272 -29 288
rect -129 238 -113 272
rect -45 238 -29 272
rect -129 200 -29 238
rect 29 272 129 288
rect 29 238 45 272
rect 113 238 129 272
rect 29 200 129 238
rect 187 272 287 288
rect 187 238 203 272
rect 271 238 287 272
rect 187 200 287 238
rect 345 272 445 288
rect 345 238 361 272
rect 429 238 445 272
rect 345 200 445 238
rect 503 272 603 288
rect 503 238 519 272
rect 587 238 603 272
rect 503 200 603 238
rect 661 272 761 288
rect 661 238 677 272
rect 745 238 761 272
rect 661 200 761 238
rect 819 272 919 288
rect 819 238 835 272
rect 903 238 919 272
rect 819 200 919 238
rect 977 272 1077 288
rect 977 238 993 272
rect 1061 238 1077 272
rect 977 200 1077 238
rect 1135 272 1235 288
rect 1135 238 1151 272
rect 1219 238 1235 272
rect 1135 200 1235 238
rect -1235 -238 -1135 -200
rect -1235 -272 -1219 -238
rect -1151 -272 -1135 -238
rect -1235 -288 -1135 -272
rect -1077 -238 -977 -200
rect -1077 -272 -1061 -238
rect -993 -272 -977 -238
rect -1077 -288 -977 -272
rect -919 -238 -819 -200
rect -919 -272 -903 -238
rect -835 -272 -819 -238
rect -919 -288 -819 -272
rect -761 -238 -661 -200
rect -761 -272 -745 -238
rect -677 -272 -661 -238
rect -761 -288 -661 -272
rect -603 -238 -503 -200
rect -603 -272 -587 -238
rect -519 -272 -503 -238
rect -603 -288 -503 -272
rect -445 -238 -345 -200
rect -445 -272 -429 -238
rect -361 -272 -345 -238
rect -445 -288 -345 -272
rect -287 -238 -187 -200
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -287 -288 -187 -272
rect -129 -238 -29 -200
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect -129 -288 -29 -272
rect 29 -238 129 -200
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 29 -288 129 -272
rect 187 -238 287 -200
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 187 -288 287 -272
rect 345 -238 445 -200
rect 345 -272 361 -238
rect 429 -272 445 -238
rect 345 -288 445 -272
rect 503 -238 603 -200
rect 503 -272 519 -238
rect 587 -272 603 -238
rect 503 -288 603 -272
rect 661 -238 761 -200
rect 661 -272 677 -238
rect 745 -272 761 -238
rect 661 -288 761 -272
rect 819 -238 919 -200
rect 819 -272 835 -238
rect 903 -272 919 -238
rect 819 -288 919 -272
rect 977 -238 1077 -200
rect 977 -272 993 -238
rect 1061 -272 1077 -238
rect 977 -288 1077 -272
rect 1135 -238 1235 -200
rect 1135 -272 1151 -238
rect 1219 -272 1235 -238
rect 1135 -288 1235 -272
<< polycont >>
rect -1219 238 -1151 272
rect -1061 238 -993 272
rect -903 238 -835 272
rect -745 238 -677 272
rect -587 238 -519 272
rect -429 238 -361 272
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect 361 238 429 272
rect 519 238 587 272
rect 677 238 745 272
rect 835 238 903 272
rect 993 238 1061 272
rect 1151 238 1219 272
rect -1219 -272 -1151 -238
rect -1061 -272 -993 -238
rect -903 -272 -835 -238
rect -745 -272 -677 -238
rect -587 -272 -519 -238
rect -429 -272 -361 -238
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
rect 361 -272 429 -238
rect 519 -272 587 -238
rect 677 -272 745 -238
rect 835 -272 903 -238
rect 993 -272 1061 -238
rect 1151 -272 1219 -238
<< locali >>
rect -1395 340 -1299 374
rect 1299 340 1395 374
rect -1395 278 -1361 340
rect 1361 278 1395 340
rect -1235 238 -1219 272
rect -1151 238 -1135 272
rect -1077 238 -1061 272
rect -993 238 -977 272
rect -919 238 -903 272
rect -835 238 -819 272
rect -761 238 -745 272
rect -677 238 -661 272
rect -603 238 -587 272
rect -519 238 -503 272
rect -445 238 -429 272
rect -361 238 -345 272
rect -287 238 -271 272
rect -203 238 -187 272
rect -129 238 -113 272
rect -45 238 -29 272
rect 29 238 45 272
rect 113 238 129 272
rect 187 238 203 272
rect 271 238 287 272
rect 345 238 361 272
rect 429 238 445 272
rect 503 238 519 272
rect 587 238 603 272
rect 661 238 677 272
rect 745 238 761 272
rect 819 238 835 272
rect 903 238 919 272
rect 977 238 993 272
rect 1061 238 1077 272
rect 1135 238 1151 272
rect 1219 238 1235 272
rect -1281 188 -1247 204
rect -1281 -204 -1247 -188
rect -1123 188 -1089 204
rect -1123 -204 -1089 -188
rect -965 188 -931 204
rect -965 -204 -931 -188
rect -807 188 -773 204
rect -807 -204 -773 -188
rect -649 188 -615 204
rect -649 -204 -615 -188
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect 615 188 649 204
rect 615 -204 649 -188
rect 773 188 807 204
rect 773 -204 807 -188
rect 931 188 965 204
rect 931 -204 965 -188
rect 1089 188 1123 204
rect 1089 -204 1123 -188
rect 1247 188 1281 204
rect 1247 -204 1281 -188
rect -1235 -272 -1219 -238
rect -1151 -272 -1135 -238
rect -1077 -272 -1061 -238
rect -993 -272 -977 -238
rect -919 -272 -903 -238
rect -835 -272 -819 -238
rect -761 -272 -745 -238
rect -677 -272 -661 -238
rect -603 -272 -587 -238
rect -519 -272 -503 -238
rect -445 -272 -429 -238
rect -361 -272 -345 -238
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 345 -272 361 -238
rect 429 -272 445 -238
rect 503 -272 519 -238
rect 587 -272 603 -238
rect 661 -272 677 -238
rect 745 -272 761 -238
rect 819 -272 835 -238
rect 903 -272 919 -238
rect 977 -272 993 -238
rect 1061 -272 1077 -238
rect 1135 -272 1151 -238
rect 1219 -272 1235 -238
rect -1395 -340 -1361 -278
rect 1361 -340 1395 -278
rect -1395 -374 -1299 -340
rect 1299 -374 1395 -340
<< viali >>
rect -1219 238 -1151 272
rect -1061 238 -993 272
rect -903 238 -835 272
rect -745 238 -677 272
rect -587 238 -519 272
rect -429 238 -361 272
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect 361 238 429 272
rect 519 238 587 272
rect 677 238 745 272
rect 835 238 903 272
rect 993 238 1061 272
rect 1151 238 1219 272
rect -1281 -188 -1247 188
rect -1123 -188 -1089 188
rect -965 -188 -931 188
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect 931 -188 965 188
rect 1089 -188 1123 188
rect 1247 -188 1281 188
rect -1219 -272 -1151 -238
rect -1061 -272 -993 -238
rect -903 -272 -835 -238
rect -745 -272 -677 -238
rect -587 -272 -519 -238
rect -429 -272 -361 -238
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
rect 361 -272 429 -238
rect 519 -272 587 -238
rect 677 -272 745 -238
rect 835 -272 903 -238
rect 993 -272 1061 -238
rect 1151 -272 1219 -238
<< metal1 >>
rect -1231 272 -1139 278
rect -1231 238 -1219 272
rect -1151 238 -1139 272
rect -1231 232 -1139 238
rect -1073 272 -981 278
rect -1073 238 -1061 272
rect -993 238 -981 272
rect -1073 232 -981 238
rect -915 272 -823 278
rect -915 238 -903 272
rect -835 238 -823 272
rect -915 232 -823 238
rect -757 272 -665 278
rect -757 238 -745 272
rect -677 238 -665 272
rect -757 232 -665 238
rect -599 272 -507 278
rect -599 238 -587 272
rect -519 238 -507 272
rect -599 232 -507 238
rect -441 272 -349 278
rect -441 238 -429 272
rect -361 238 -349 272
rect -441 232 -349 238
rect -283 272 -191 278
rect -283 238 -271 272
rect -203 238 -191 272
rect -283 232 -191 238
rect -125 272 -33 278
rect -125 238 -113 272
rect -45 238 -33 272
rect -125 232 -33 238
rect 33 272 125 278
rect 33 238 45 272
rect 113 238 125 272
rect 33 232 125 238
rect 191 272 283 278
rect 191 238 203 272
rect 271 238 283 272
rect 191 232 283 238
rect 349 272 441 278
rect 349 238 361 272
rect 429 238 441 272
rect 349 232 441 238
rect 507 272 599 278
rect 507 238 519 272
rect 587 238 599 272
rect 507 232 599 238
rect 665 272 757 278
rect 665 238 677 272
rect 745 238 757 272
rect 665 232 757 238
rect 823 272 915 278
rect 823 238 835 272
rect 903 238 915 272
rect 823 232 915 238
rect 981 272 1073 278
rect 981 238 993 272
rect 1061 238 1073 272
rect 981 232 1073 238
rect 1139 272 1231 278
rect 1139 238 1151 272
rect 1219 238 1231 272
rect 1139 232 1231 238
rect -1287 188 -1241 200
rect -1287 -188 -1281 188
rect -1247 -188 -1241 188
rect -1287 -200 -1241 -188
rect -1129 188 -1083 200
rect -1129 -188 -1123 188
rect -1089 -188 -1083 188
rect -1129 -200 -1083 -188
rect -971 188 -925 200
rect -971 -188 -965 188
rect -931 -188 -925 188
rect -971 -200 -925 -188
rect -813 188 -767 200
rect -813 -188 -807 188
rect -773 -188 -767 188
rect -813 -200 -767 -188
rect -655 188 -609 200
rect -655 -188 -649 188
rect -615 -188 -609 188
rect -655 -200 -609 -188
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect 609 188 655 200
rect 609 -188 615 188
rect 649 -188 655 188
rect 609 -200 655 -188
rect 767 188 813 200
rect 767 -188 773 188
rect 807 -188 813 188
rect 767 -200 813 -188
rect 925 188 971 200
rect 925 -188 931 188
rect 965 -188 971 188
rect 925 -200 971 -188
rect 1083 188 1129 200
rect 1083 -188 1089 188
rect 1123 -188 1129 188
rect 1083 -200 1129 -188
rect 1241 188 1287 200
rect 1241 -188 1247 188
rect 1281 -188 1287 188
rect 1241 -200 1287 -188
rect -1231 -238 -1139 -232
rect -1231 -272 -1219 -238
rect -1151 -272 -1139 -238
rect -1231 -278 -1139 -272
rect -1073 -238 -981 -232
rect -1073 -272 -1061 -238
rect -993 -272 -981 -238
rect -1073 -278 -981 -272
rect -915 -238 -823 -232
rect -915 -272 -903 -238
rect -835 -272 -823 -238
rect -915 -278 -823 -272
rect -757 -238 -665 -232
rect -757 -272 -745 -238
rect -677 -272 -665 -238
rect -757 -278 -665 -272
rect -599 -238 -507 -232
rect -599 -272 -587 -238
rect -519 -272 -507 -238
rect -599 -278 -507 -272
rect -441 -238 -349 -232
rect -441 -272 -429 -238
rect -361 -272 -349 -238
rect -441 -278 -349 -272
rect -283 -238 -191 -232
rect -283 -272 -271 -238
rect -203 -272 -191 -238
rect -283 -278 -191 -272
rect -125 -238 -33 -232
rect -125 -272 -113 -238
rect -45 -272 -33 -238
rect -125 -278 -33 -272
rect 33 -238 125 -232
rect 33 -272 45 -238
rect 113 -272 125 -238
rect 33 -278 125 -272
rect 191 -238 283 -232
rect 191 -272 203 -238
rect 271 -272 283 -238
rect 191 -278 283 -272
rect 349 -238 441 -232
rect 349 -272 361 -238
rect 429 -272 441 -238
rect 349 -278 441 -272
rect 507 -238 599 -232
rect 507 -272 519 -238
rect 587 -272 599 -238
rect 507 -278 599 -272
rect 665 -238 757 -232
rect 665 -272 677 -238
rect 745 -272 757 -238
rect 665 -278 757 -272
rect 823 -238 915 -232
rect 823 -272 835 -238
rect 903 -272 915 -238
rect 823 -278 915 -272
rect 981 -238 1073 -232
rect 981 -272 993 -238
rect 1061 -272 1073 -238
rect 981 -278 1073 -272
rect 1139 -238 1231 -232
rect 1139 -272 1151 -238
rect 1219 -272 1231 -238
rect 1139 -278 1231 -272
<< properties >>
string FIXED_BBOX -1378 -357 1378 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.5 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
