magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< pwell >>
rect 890 900 1436 906
rect 890 850 1480 900
rect 890 840 1436 850
rect 890 390 1436 396
rect 890 340 1474 390
rect 890 330 1436 340
<< poly >>
rect 890 890 1436 906
rect 890 856 906 890
rect 940 856 1098 890
rect 1132 856 1290 890
rect 1324 856 1436 890
rect 890 840 1436 856
rect 890 380 1436 396
rect 890 346 1002 380
rect 1036 346 1194 380
rect 1228 346 1386 380
rect 1420 346 1436 380
rect 890 330 1436 346
<< polycont >>
rect 906 856 940 890
rect 1098 856 1132 890
rect 1290 856 1324 890
rect 1002 346 1036 380
rect 1194 346 1228 380
rect 1386 346 1420 380
<< locali >>
rect 890 856 906 890
rect 940 856 1098 890
rect 1132 856 1290 890
rect 1324 856 1436 890
rect 890 346 1002 380
rect 1036 346 1194 380
rect 1228 346 1386 380
rect 1420 346 1436 380
<< viali >>
rect 906 856 940 890
rect 1098 856 1132 890
rect 1290 856 1324 890
rect 1002 346 1036 380
rect 1194 346 1228 380
rect 1386 346 1420 380
<< metal1 >>
rect 760 890 1570 900
rect 760 856 906 890
rect 940 856 1098 890
rect 1132 856 1290 890
rect 1324 856 1570 890
rect 760 850 1570 856
rect 760 390 810 850
rect 934 642 944 818
rect 998 642 1008 818
rect 1126 642 1136 818
rect 1190 642 1200 818
rect 1318 642 1328 818
rect 1382 642 1392 818
rect 838 418 848 594
rect 902 418 912 594
rect 1030 418 1040 594
rect 1094 418 1104 594
rect 1222 418 1232 594
rect 1286 418 1296 594
rect 1414 418 1424 594
rect 1478 418 1488 594
rect 1520 390 1570 850
rect 760 380 1570 390
rect 760 346 1002 380
rect 1036 346 1194 380
rect 1228 346 1386 380
rect 1420 346 1570 380
rect 760 340 1570 346
<< via1 >>
rect 944 642 998 818
rect 1136 642 1190 818
rect 1328 642 1382 818
rect 848 418 902 594
rect 1040 418 1094 594
rect 1232 418 1286 594
rect 1424 418 1478 594
<< metal2 >>
rect 944 818 998 828
rect 944 632 998 642
rect 1136 818 1190 828
rect 1136 632 1190 642
rect 1328 818 1382 828
rect 1328 632 1382 642
rect 848 594 902 604
rect 848 408 902 418
rect 1040 594 1094 604
rect 1040 408 1094 418
rect 1232 594 1286 604
rect 1232 408 1286 418
rect 1424 594 1478 604
rect 1424 408 1478 418
use sky130_fd_pr__nfet_01v8_lvt_V6SMGN  sky130_fd_pr__nfet_01v8_lvt_V6SMGN_0
timestamp 1654768133
transform 1 0 1163 0 1 618
box -455 -410 455 410
<< end >>
