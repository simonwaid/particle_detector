magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< metal4 >>
rect -3351 1559 3351 1600
rect -3351 -1559 3095 1559
rect 3331 -1559 3351 1559
rect -3351 -1600 3351 -1559
<< via4 >>
rect 3095 -1559 3331 1559
<< mimcap2 >>
rect -3251 1460 2749 1500
rect -3251 -1460 -3211 1460
rect 2709 -1460 2749 1460
rect -3251 -1500 2749 -1460
<< mimcap2contact >>
rect -3211 -1460 2709 1460
<< metal5 >>
rect 3053 1559 3373 1601
rect -3235 1460 2733 1484
rect -3235 -1460 -3211 1460
rect 2709 -1460 2733 1460
rect -3235 -1484 2733 -1460
rect 3053 -1559 3095 1559
rect 3331 -1559 3373 1559
rect 3053 -1601 3373 -1559
<< properties >>
string FIXED_BBOX -3351 -1600 2849 1600
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 15 val 917.1 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
