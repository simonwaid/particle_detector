magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< error_p >>
rect -1150 272 -1092 278
rect -1032 272 -974 278
rect -914 272 -856 278
rect -796 272 -738 278
rect -678 272 -620 278
rect -560 272 -502 278
rect -442 272 -384 278
rect -324 272 -266 278
rect -206 272 -148 278
rect -88 272 -30 278
rect 30 272 88 278
rect 148 272 206 278
rect 266 272 324 278
rect 384 272 442 278
rect 502 272 560 278
rect 620 272 678 278
rect 738 272 796 278
rect 856 272 914 278
rect 974 272 1032 278
rect 1092 272 1150 278
rect -1150 238 -1138 272
rect -1032 238 -1020 272
rect -914 238 -902 272
rect -796 238 -784 272
rect -678 238 -666 272
rect -560 238 -548 272
rect -442 238 -430 272
rect -324 238 -312 272
rect -206 238 -194 272
rect -88 238 -76 272
rect 30 238 42 272
rect 148 238 160 272
rect 266 238 278 272
rect 384 238 396 272
rect 502 238 514 272
rect 620 238 632 272
rect 738 238 750 272
rect 856 238 868 272
rect 974 238 986 272
rect 1092 238 1104 272
rect -1150 232 -1092 238
rect -1032 232 -974 238
rect -914 232 -856 238
rect -796 232 -738 238
rect -678 232 -620 238
rect -560 232 -502 238
rect -442 232 -384 238
rect -324 232 -266 238
rect -206 232 -148 238
rect -88 232 -30 238
rect 30 232 88 238
rect 148 232 206 238
rect 266 232 324 238
rect 384 232 442 238
rect 502 232 560 238
rect 620 232 678 238
rect 738 232 796 238
rect 856 232 914 238
rect 974 232 1032 238
rect 1092 232 1150 238
rect -1150 -238 -1092 -232
rect -1032 -238 -974 -232
rect -914 -238 -856 -232
rect -796 -238 -738 -232
rect -678 -238 -620 -232
rect -560 -238 -502 -232
rect -442 -238 -384 -232
rect -324 -238 -266 -232
rect -206 -238 -148 -232
rect -88 -238 -30 -232
rect 30 -238 88 -232
rect 148 -238 206 -232
rect 266 -238 324 -232
rect 384 -238 442 -232
rect 502 -238 560 -232
rect 620 -238 678 -232
rect 738 -238 796 -232
rect 856 -238 914 -232
rect 974 -238 1032 -232
rect 1092 -238 1150 -232
rect -1150 -272 -1138 -238
rect -1032 -272 -1020 -238
rect -914 -272 -902 -238
rect -796 -272 -784 -238
rect -678 -272 -666 -238
rect -560 -272 -548 -238
rect -442 -272 -430 -238
rect -324 -272 -312 -238
rect -206 -272 -194 -238
rect -88 -272 -76 -238
rect 30 -272 42 -238
rect 148 -272 160 -238
rect 266 -272 278 -238
rect 384 -272 396 -238
rect 502 -272 514 -238
rect 620 -272 632 -238
rect 738 -272 750 -238
rect 856 -272 868 -238
rect 974 -272 986 -238
rect 1092 -272 1104 -238
rect -1150 -278 -1092 -272
rect -1032 -278 -974 -272
rect -914 -278 -856 -272
rect -796 -278 -738 -272
rect -678 -278 -620 -272
rect -560 -278 -502 -272
rect -442 -278 -384 -272
rect -324 -278 -266 -272
rect -206 -278 -148 -272
rect -88 -278 -30 -272
rect 30 -278 88 -272
rect 148 -278 206 -272
rect 266 -278 324 -272
rect 384 -278 442 -272
rect 502 -278 560 -272
rect 620 -278 678 -272
rect 738 -278 796 -272
rect 856 -278 914 -272
rect 974 -278 1032 -272
rect 1092 -278 1150 -272
<< pwell >>
rect -1347 -410 1347 410
<< nmos >>
rect -1151 -200 -1091 200
rect -1033 -200 -973 200
rect -915 -200 -855 200
rect -797 -200 -737 200
rect -679 -200 -619 200
rect -561 -200 -501 200
rect -443 -200 -383 200
rect -325 -200 -265 200
rect -207 -200 -147 200
rect -89 -200 -29 200
rect 29 -200 89 200
rect 147 -200 207 200
rect 265 -200 325 200
rect 383 -200 443 200
rect 501 -200 561 200
rect 619 -200 679 200
rect 737 -200 797 200
rect 855 -200 915 200
rect 973 -200 1033 200
rect 1091 -200 1151 200
<< ndiff >>
rect -1209 188 -1151 200
rect -1209 -188 -1197 188
rect -1163 -188 -1151 188
rect -1209 -200 -1151 -188
rect -1091 188 -1033 200
rect -1091 -188 -1079 188
rect -1045 -188 -1033 188
rect -1091 -200 -1033 -188
rect -973 188 -915 200
rect -973 -188 -961 188
rect -927 -188 -915 188
rect -973 -200 -915 -188
rect -855 188 -797 200
rect -855 -188 -843 188
rect -809 -188 -797 188
rect -855 -200 -797 -188
rect -737 188 -679 200
rect -737 -188 -725 188
rect -691 -188 -679 188
rect -737 -200 -679 -188
rect -619 188 -561 200
rect -619 -188 -607 188
rect -573 -188 -561 188
rect -619 -200 -561 -188
rect -501 188 -443 200
rect -501 -188 -489 188
rect -455 -188 -443 188
rect -501 -200 -443 -188
rect -383 188 -325 200
rect -383 -188 -371 188
rect -337 -188 -325 188
rect -383 -200 -325 -188
rect -265 188 -207 200
rect -265 -188 -253 188
rect -219 -188 -207 188
rect -265 -200 -207 -188
rect -147 188 -89 200
rect -147 -188 -135 188
rect -101 -188 -89 188
rect -147 -200 -89 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 89 188 147 200
rect 89 -188 101 188
rect 135 -188 147 188
rect 89 -200 147 -188
rect 207 188 265 200
rect 207 -188 219 188
rect 253 -188 265 188
rect 207 -200 265 -188
rect 325 188 383 200
rect 325 -188 337 188
rect 371 -188 383 188
rect 325 -200 383 -188
rect 443 188 501 200
rect 443 -188 455 188
rect 489 -188 501 188
rect 443 -200 501 -188
rect 561 188 619 200
rect 561 -188 573 188
rect 607 -188 619 188
rect 561 -200 619 -188
rect 679 188 737 200
rect 679 -188 691 188
rect 725 -188 737 188
rect 679 -200 737 -188
rect 797 188 855 200
rect 797 -188 809 188
rect 843 -188 855 188
rect 797 -200 855 -188
rect 915 188 973 200
rect 915 -188 927 188
rect 961 -188 973 188
rect 915 -200 973 -188
rect 1033 188 1091 200
rect 1033 -188 1045 188
rect 1079 -188 1091 188
rect 1033 -200 1091 -188
rect 1151 188 1209 200
rect 1151 -188 1163 188
rect 1197 -188 1209 188
rect 1151 -200 1209 -188
<< ndiffc >>
rect -1197 -188 -1163 188
rect -1079 -188 -1045 188
rect -961 -188 -927 188
rect -843 -188 -809 188
rect -725 -188 -691 188
rect -607 -188 -573 188
rect -489 -188 -455 188
rect -371 -188 -337 188
rect -253 -188 -219 188
rect -135 -188 -101 188
rect -17 -188 17 188
rect 101 -188 135 188
rect 219 -188 253 188
rect 337 -188 371 188
rect 455 -188 489 188
rect 573 -188 607 188
rect 691 -188 725 188
rect 809 -188 843 188
rect 927 -188 961 188
rect 1045 -188 1079 188
rect 1163 -188 1197 188
<< psubdiff >>
rect -1311 340 -1215 374
rect 1215 340 1311 374
rect -1311 278 -1277 340
rect 1277 278 1311 340
rect -1311 -340 -1277 -278
rect 1277 -340 1311 -278
rect -1311 -374 -1215 -340
rect 1215 -374 1311 -340
<< psubdiffcont >>
rect -1215 340 1215 374
rect -1311 -278 -1277 278
rect 1277 -278 1311 278
rect -1215 -374 1215 -340
<< poly >>
rect -1154 272 -1088 288
rect -1154 238 -1138 272
rect -1104 238 -1088 272
rect -1154 222 -1088 238
rect -1036 272 -970 288
rect -1036 238 -1020 272
rect -986 238 -970 272
rect -1036 222 -970 238
rect -918 272 -852 288
rect -918 238 -902 272
rect -868 238 -852 272
rect -918 222 -852 238
rect -800 272 -734 288
rect -800 238 -784 272
rect -750 238 -734 272
rect -800 222 -734 238
rect -682 272 -616 288
rect -682 238 -666 272
rect -632 238 -616 272
rect -682 222 -616 238
rect -564 272 -498 288
rect -564 238 -548 272
rect -514 238 -498 272
rect -564 222 -498 238
rect -446 272 -380 288
rect -446 238 -430 272
rect -396 238 -380 272
rect -446 222 -380 238
rect -328 272 -262 288
rect -328 238 -312 272
rect -278 238 -262 272
rect -328 222 -262 238
rect -210 272 -144 288
rect -210 238 -194 272
rect -160 238 -144 272
rect -210 222 -144 238
rect -92 272 -26 288
rect -92 238 -76 272
rect -42 238 -26 272
rect -92 222 -26 238
rect 26 272 92 288
rect 26 238 42 272
rect 76 238 92 272
rect 26 222 92 238
rect 144 272 210 288
rect 144 238 160 272
rect 194 238 210 272
rect 144 222 210 238
rect 262 272 328 288
rect 262 238 278 272
rect 312 238 328 272
rect 262 222 328 238
rect 380 272 446 288
rect 380 238 396 272
rect 430 238 446 272
rect 380 222 446 238
rect 498 272 564 288
rect 498 238 514 272
rect 548 238 564 272
rect 498 222 564 238
rect 616 272 682 288
rect 616 238 632 272
rect 666 238 682 272
rect 616 222 682 238
rect 734 272 800 288
rect 734 238 750 272
rect 784 238 800 272
rect 734 222 800 238
rect 852 272 918 288
rect 852 238 868 272
rect 902 238 918 272
rect 852 222 918 238
rect 970 272 1036 288
rect 970 238 986 272
rect 1020 238 1036 272
rect 970 222 1036 238
rect 1088 272 1154 288
rect 1088 238 1104 272
rect 1138 238 1154 272
rect 1088 222 1154 238
rect -1151 200 -1091 222
rect -1033 200 -973 222
rect -915 200 -855 222
rect -797 200 -737 222
rect -679 200 -619 222
rect -561 200 -501 222
rect -443 200 -383 222
rect -325 200 -265 222
rect -207 200 -147 222
rect -89 200 -29 222
rect 29 200 89 222
rect 147 200 207 222
rect 265 200 325 222
rect 383 200 443 222
rect 501 200 561 222
rect 619 200 679 222
rect 737 200 797 222
rect 855 200 915 222
rect 973 200 1033 222
rect 1091 200 1151 222
rect -1151 -222 -1091 -200
rect -1033 -222 -973 -200
rect -915 -222 -855 -200
rect -797 -222 -737 -200
rect -679 -222 -619 -200
rect -561 -222 -501 -200
rect -443 -222 -383 -200
rect -325 -222 -265 -200
rect -207 -222 -147 -200
rect -89 -222 -29 -200
rect 29 -222 89 -200
rect 147 -222 207 -200
rect 265 -222 325 -200
rect 383 -222 443 -200
rect 501 -222 561 -200
rect 619 -222 679 -200
rect 737 -222 797 -200
rect 855 -222 915 -200
rect 973 -222 1033 -200
rect 1091 -222 1151 -200
rect -1154 -238 -1088 -222
rect -1154 -272 -1138 -238
rect -1104 -272 -1088 -238
rect -1154 -288 -1088 -272
rect -1036 -238 -970 -222
rect -1036 -272 -1020 -238
rect -986 -272 -970 -238
rect -1036 -288 -970 -272
rect -918 -238 -852 -222
rect -918 -272 -902 -238
rect -868 -272 -852 -238
rect -918 -288 -852 -272
rect -800 -238 -734 -222
rect -800 -272 -784 -238
rect -750 -272 -734 -238
rect -800 -288 -734 -272
rect -682 -238 -616 -222
rect -682 -272 -666 -238
rect -632 -272 -616 -238
rect -682 -288 -616 -272
rect -564 -238 -498 -222
rect -564 -272 -548 -238
rect -514 -272 -498 -238
rect -564 -288 -498 -272
rect -446 -238 -380 -222
rect -446 -272 -430 -238
rect -396 -272 -380 -238
rect -446 -288 -380 -272
rect -328 -238 -262 -222
rect -328 -272 -312 -238
rect -278 -272 -262 -238
rect -328 -288 -262 -272
rect -210 -238 -144 -222
rect -210 -272 -194 -238
rect -160 -272 -144 -238
rect -210 -288 -144 -272
rect -92 -238 -26 -222
rect -92 -272 -76 -238
rect -42 -272 -26 -238
rect -92 -288 -26 -272
rect 26 -238 92 -222
rect 26 -272 42 -238
rect 76 -272 92 -238
rect 26 -288 92 -272
rect 144 -238 210 -222
rect 144 -272 160 -238
rect 194 -272 210 -238
rect 144 -288 210 -272
rect 262 -238 328 -222
rect 262 -272 278 -238
rect 312 -272 328 -238
rect 262 -288 328 -272
rect 380 -238 446 -222
rect 380 -272 396 -238
rect 430 -272 446 -238
rect 380 -288 446 -272
rect 498 -238 564 -222
rect 498 -272 514 -238
rect 548 -272 564 -238
rect 498 -288 564 -272
rect 616 -238 682 -222
rect 616 -272 632 -238
rect 666 -272 682 -238
rect 616 -288 682 -272
rect 734 -238 800 -222
rect 734 -272 750 -238
rect 784 -272 800 -238
rect 734 -288 800 -272
rect 852 -238 918 -222
rect 852 -272 868 -238
rect 902 -272 918 -238
rect 852 -288 918 -272
rect 970 -238 1036 -222
rect 970 -272 986 -238
rect 1020 -272 1036 -238
rect 970 -288 1036 -272
rect 1088 -238 1154 -222
rect 1088 -272 1104 -238
rect 1138 -272 1154 -238
rect 1088 -288 1154 -272
<< polycont >>
rect -1138 238 -1104 272
rect -1020 238 -986 272
rect -902 238 -868 272
rect -784 238 -750 272
rect -666 238 -632 272
rect -548 238 -514 272
rect -430 238 -396 272
rect -312 238 -278 272
rect -194 238 -160 272
rect -76 238 -42 272
rect 42 238 76 272
rect 160 238 194 272
rect 278 238 312 272
rect 396 238 430 272
rect 514 238 548 272
rect 632 238 666 272
rect 750 238 784 272
rect 868 238 902 272
rect 986 238 1020 272
rect 1104 238 1138 272
rect -1138 -272 -1104 -238
rect -1020 -272 -986 -238
rect -902 -272 -868 -238
rect -784 -272 -750 -238
rect -666 -272 -632 -238
rect -548 -272 -514 -238
rect -430 -272 -396 -238
rect -312 -272 -278 -238
rect -194 -272 -160 -238
rect -76 -272 -42 -238
rect 42 -272 76 -238
rect 160 -272 194 -238
rect 278 -272 312 -238
rect 396 -272 430 -238
rect 514 -272 548 -238
rect 632 -272 666 -238
rect 750 -272 784 -238
rect 868 -272 902 -238
rect 986 -272 1020 -238
rect 1104 -272 1138 -238
<< locali >>
rect -1311 340 -1215 374
rect 1215 340 1311 374
rect -1311 278 -1277 340
rect 1277 278 1311 340
rect -1154 238 -1138 272
rect -1104 238 -1088 272
rect -1036 238 -1020 272
rect -986 238 -970 272
rect -918 238 -902 272
rect -868 238 -852 272
rect -800 238 -784 272
rect -750 238 -734 272
rect -682 238 -666 272
rect -632 238 -616 272
rect -564 238 -548 272
rect -514 238 -498 272
rect -446 238 -430 272
rect -396 238 -380 272
rect -328 238 -312 272
rect -278 238 -262 272
rect -210 238 -194 272
rect -160 238 -144 272
rect -92 238 -76 272
rect -42 238 -26 272
rect 26 238 42 272
rect 76 238 92 272
rect 144 238 160 272
rect 194 238 210 272
rect 262 238 278 272
rect 312 238 328 272
rect 380 238 396 272
rect 430 238 446 272
rect 498 238 514 272
rect 548 238 564 272
rect 616 238 632 272
rect 666 238 682 272
rect 734 238 750 272
rect 784 238 800 272
rect 852 238 868 272
rect 902 238 918 272
rect 970 238 986 272
rect 1020 238 1036 272
rect 1088 238 1104 272
rect 1138 238 1154 272
rect -1197 188 -1163 204
rect -1197 -204 -1163 -188
rect -1079 188 -1045 204
rect -1079 -204 -1045 -188
rect -961 188 -927 204
rect -961 -204 -927 -188
rect -843 188 -809 204
rect -843 -204 -809 -188
rect -725 188 -691 204
rect -725 -204 -691 -188
rect -607 188 -573 204
rect -607 -204 -573 -188
rect -489 188 -455 204
rect -489 -204 -455 -188
rect -371 188 -337 204
rect -371 -204 -337 -188
rect -253 188 -219 204
rect -253 -204 -219 -188
rect -135 188 -101 204
rect -135 -204 -101 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 101 188 135 204
rect 101 -204 135 -188
rect 219 188 253 204
rect 219 -204 253 -188
rect 337 188 371 204
rect 337 -204 371 -188
rect 455 188 489 204
rect 455 -204 489 -188
rect 573 188 607 204
rect 573 -204 607 -188
rect 691 188 725 204
rect 691 -204 725 -188
rect 809 188 843 204
rect 809 -204 843 -188
rect 927 188 961 204
rect 927 -204 961 -188
rect 1045 188 1079 204
rect 1045 -204 1079 -188
rect 1163 188 1197 204
rect 1163 -204 1197 -188
rect -1154 -272 -1138 -238
rect -1104 -272 -1088 -238
rect -1036 -272 -1020 -238
rect -986 -272 -970 -238
rect -918 -272 -902 -238
rect -868 -272 -852 -238
rect -800 -272 -784 -238
rect -750 -272 -734 -238
rect -682 -272 -666 -238
rect -632 -272 -616 -238
rect -564 -272 -548 -238
rect -514 -272 -498 -238
rect -446 -272 -430 -238
rect -396 -272 -380 -238
rect -328 -272 -312 -238
rect -278 -272 -262 -238
rect -210 -272 -194 -238
rect -160 -272 -144 -238
rect -92 -272 -76 -238
rect -42 -272 -26 -238
rect 26 -272 42 -238
rect 76 -272 92 -238
rect 144 -272 160 -238
rect 194 -272 210 -238
rect 262 -272 278 -238
rect 312 -272 328 -238
rect 380 -272 396 -238
rect 430 -272 446 -238
rect 498 -272 514 -238
rect 548 -272 564 -238
rect 616 -272 632 -238
rect 666 -272 682 -238
rect 734 -272 750 -238
rect 784 -272 800 -238
rect 852 -272 868 -238
rect 902 -272 918 -238
rect 970 -272 986 -238
rect 1020 -272 1036 -238
rect 1088 -272 1104 -238
rect 1138 -272 1154 -238
rect -1311 -340 -1277 -278
rect 1277 -340 1311 -278
rect -1311 -374 -1215 -340
rect 1215 -374 1311 -340
<< viali >>
rect -1138 238 -1104 272
rect -1020 238 -986 272
rect -902 238 -868 272
rect -784 238 -750 272
rect -666 238 -632 272
rect -548 238 -514 272
rect -430 238 -396 272
rect -312 238 -278 272
rect -194 238 -160 272
rect -76 238 -42 272
rect 42 238 76 272
rect 160 238 194 272
rect 278 238 312 272
rect 396 238 430 272
rect 514 238 548 272
rect 632 238 666 272
rect 750 238 784 272
rect 868 238 902 272
rect 986 238 1020 272
rect 1104 238 1138 272
rect -1197 -188 -1163 188
rect -1079 -188 -1045 188
rect -961 -188 -927 188
rect -843 -188 -809 188
rect -725 -188 -691 188
rect -607 -188 -573 188
rect -489 -188 -455 188
rect -371 -188 -337 188
rect -253 -188 -219 188
rect -135 -188 -101 188
rect -17 -188 17 188
rect 101 -188 135 188
rect 219 -188 253 188
rect 337 -188 371 188
rect 455 -188 489 188
rect 573 -188 607 188
rect 691 -188 725 188
rect 809 -188 843 188
rect 927 -188 961 188
rect 1045 -188 1079 188
rect 1163 -188 1197 188
rect -1138 -272 -1104 -238
rect -1020 -272 -986 -238
rect -902 -272 -868 -238
rect -784 -272 -750 -238
rect -666 -272 -632 -238
rect -548 -272 -514 -238
rect -430 -272 -396 -238
rect -312 -272 -278 -238
rect -194 -272 -160 -238
rect -76 -272 -42 -238
rect 42 -272 76 -238
rect 160 -272 194 -238
rect 278 -272 312 -238
rect 396 -272 430 -238
rect 514 -272 548 -238
rect 632 -272 666 -238
rect 750 -272 784 -238
rect 868 -272 902 -238
rect 986 -272 1020 -238
rect 1104 -272 1138 -238
<< metal1 >>
rect -1150 272 -1092 278
rect -1150 238 -1138 272
rect -1104 238 -1092 272
rect -1150 232 -1092 238
rect -1032 272 -974 278
rect -1032 238 -1020 272
rect -986 238 -974 272
rect -1032 232 -974 238
rect -914 272 -856 278
rect -914 238 -902 272
rect -868 238 -856 272
rect -914 232 -856 238
rect -796 272 -738 278
rect -796 238 -784 272
rect -750 238 -738 272
rect -796 232 -738 238
rect -678 272 -620 278
rect -678 238 -666 272
rect -632 238 -620 272
rect -678 232 -620 238
rect -560 272 -502 278
rect -560 238 -548 272
rect -514 238 -502 272
rect -560 232 -502 238
rect -442 272 -384 278
rect -442 238 -430 272
rect -396 238 -384 272
rect -442 232 -384 238
rect -324 272 -266 278
rect -324 238 -312 272
rect -278 238 -266 272
rect -324 232 -266 238
rect -206 272 -148 278
rect -206 238 -194 272
rect -160 238 -148 272
rect -206 232 -148 238
rect -88 272 -30 278
rect -88 238 -76 272
rect -42 238 -30 272
rect -88 232 -30 238
rect 30 272 88 278
rect 30 238 42 272
rect 76 238 88 272
rect 30 232 88 238
rect 148 272 206 278
rect 148 238 160 272
rect 194 238 206 272
rect 148 232 206 238
rect 266 272 324 278
rect 266 238 278 272
rect 312 238 324 272
rect 266 232 324 238
rect 384 272 442 278
rect 384 238 396 272
rect 430 238 442 272
rect 384 232 442 238
rect 502 272 560 278
rect 502 238 514 272
rect 548 238 560 272
rect 502 232 560 238
rect 620 272 678 278
rect 620 238 632 272
rect 666 238 678 272
rect 620 232 678 238
rect 738 272 796 278
rect 738 238 750 272
rect 784 238 796 272
rect 738 232 796 238
rect 856 272 914 278
rect 856 238 868 272
rect 902 238 914 272
rect 856 232 914 238
rect 974 272 1032 278
rect 974 238 986 272
rect 1020 238 1032 272
rect 974 232 1032 238
rect 1092 272 1150 278
rect 1092 238 1104 272
rect 1138 238 1150 272
rect 1092 232 1150 238
rect -1203 188 -1157 200
rect -1203 -188 -1197 188
rect -1163 -188 -1157 188
rect -1203 -200 -1157 -188
rect -1085 188 -1039 200
rect -1085 -188 -1079 188
rect -1045 -188 -1039 188
rect -1085 -200 -1039 -188
rect -967 188 -921 200
rect -967 -188 -961 188
rect -927 -188 -921 188
rect -967 -200 -921 -188
rect -849 188 -803 200
rect -849 -188 -843 188
rect -809 -188 -803 188
rect -849 -200 -803 -188
rect -731 188 -685 200
rect -731 -188 -725 188
rect -691 -188 -685 188
rect -731 -200 -685 -188
rect -613 188 -567 200
rect -613 -188 -607 188
rect -573 -188 -567 188
rect -613 -200 -567 -188
rect -495 188 -449 200
rect -495 -188 -489 188
rect -455 -188 -449 188
rect -495 -200 -449 -188
rect -377 188 -331 200
rect -377 -188 -371 188
rect -337 -188 -331 188
rect -377 -200 -331 -188
rect -259 188 -213 200
rect -259 -188 -253 188
rect -219 -188 -213 188
rect -259 -200 -213 -188
rect -141 188 -95 200
rect -141 -188 -135 188
rect -101 -188 -95 188
rect -141 -200 -95 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 95 188 141 200
rect 95 -188 101 188
rect 135 -188 141 188
rect 95 -200 141 -188
rect 213 188 259 200
rect 213 -188 219 188
rect 253 -188 259 188
rect 213 -200 259 -188
rect 331 188 377 200
rect 331 -188 337 188
rect 371 -188 377 188
rect 331 -200 377 -188
rect 449 188 495 200
rect 449 -188 455 188
rect 489 -188 495 188
rect 449 -200 495 -188
rect 567 188 613 200
rect 567 -188 573 188
rect 607 -188 613 188
rect 567 -200 613 -188
rect 685 188 731 200
rect 685 -188 691 188
rect 725 -188 731 188
rect 685 -200 731 -188
rect 803 188 849 200
rect 803 -188 809 188
rect 843 -188 849 188
rect 803 -200 849 -188
rect 921 188 967 200
rect 921 -188 927 188
rect 961 -188 967 188
rect 921 -200 967 -188
rect 1039 188 1085 200
rect 1039 -188 1045 188
rect 1079 -188 1085 188
rect 1039 -200 1085 -188
rect 1157 188 1203 200
rect 1157 -188 1163 188
rect 1197 -188 1203 188
rect 1157 -200 1203 -188
rect -1150 -238 -1092 -232
rect -1150 -272 -1138 -238
rect -1104 -272 -1092 -238
rect -1150 -278 -1092 -272
rect -1032 -238 -974 -232
rect -1032 -272 -1020 -238
rect -986 -272 -974 -238
rect -1032 -278 -974 -272
rect -914 -238 -856 -232
rect -914 -272 -902 -238
rect -868 -272 -856 -238
rect -914 -278 -856 -272
rect -796 -238 -738 -232
rect -796 -272 -784 -238
rect -750 -272 -738 -238
rect -796 -278 -738 -272
rect -678 -238 -620 -232
rect -678 -272 -666 -238
rect -632 -272 -620 -238
rect -678 -278 -620 -272
rect -560 -238 -502 -232
rect -560 -272 -548 -238
rect -514 -272 -502 -238
rect -560 -278 -502 -272
rect -442 -238 -384 -232
rect -442 -272 -430 -238
rect -396 -272 -384 -238
rect -442 -278 -384 -272
rect -324 -238 -266 -232
rect -324 -272 -312 -238
rect -278 -272 -266 -238
rect -324 -278 -266 -272
rect -206 -238 -148 -232
rect -206 -272 -194 -238
rect -160 -272 -148 -238
rect -206 -278 -148 -272
rect -88 -238 -30 -232
rect -88 -272 -76 -238
rect -42 -272 -30 -238
rect -88 -278 -30 -272
rect 30 -238 88 -232
rect 30 -272 42 -238
rect 76 -272 88 -238
rect 30 -278 88 -272
rect 148 -238 206 -232
rect 148 -272 160 -238
rect 194 -272 206 -238
rect 148 -278 206 -272
rect 266 -238 324 -232
rect 266 -272 278 -238
rect 312 -272 324 -238
rect 266 -278 324 -272
rect 384 -238 442 -232
rect 384 -272 396 -238
rect 430 -272 442 -238
rect 384 -278 442 -272
rect 502 -238 560 -232
rect 502 -272 514 -238
rect 548 -272 560 -238
rect 502 -278 560 -272
rect 620 -238 678 -232
rect 620 -272 632 -238
rect 666 -272 678 -238
rect 620 -278 678 -272
rect 738 -238 796 -232
rect 738 -272 750 -238
rect 784 -272 796 -238
rect 738 -278 796 -272
rect 856 -238 914 -232
rect 856 -272 868 -238
rect 902 -272 914 -238
rect 856 -278 914 -272
rect 974 -238 1032 -232
rect 974 -272 986 -238
rect 1020 -272 1032 -238
rect 974 -278 1032 -272
rect 1092 -238 1150 -232
rect 1092 -272 1104 -238
rect 1138 -272 1150 -238
rect 1092 -278 1150 -272
<< properties >>
string FIXED_BBOX -1294 -357 1294 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.3 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
