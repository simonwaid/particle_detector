* SPICE3 file created from outd_stage2.ext - technology: sky130A

X0 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X7 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X8 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X9 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X10 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X11 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X12 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X13 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X14 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X15 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X16 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X39 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X40 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X41 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X42 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X43 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X45 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X48 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X51 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X53 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X56 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X57 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X58 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X59 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X61 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X64 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X65 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X66 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X67 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X69 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X70 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X72 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X75 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X76 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X77 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X80 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X83 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X85 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X90 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X92 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X93 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X94 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X98 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X99 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X100 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X101 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X102 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X104 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X105 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X106 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X107 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X108 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X109 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X110 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X111 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X112 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X113 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X114 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X115 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X116 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X117 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X118 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X119 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X120 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X121 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X122 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X123 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X124 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X125 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X126 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X127 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X128 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X129 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X130 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X131 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X132 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X133 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X134 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X135 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X136 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X137 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X138 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X139 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X140 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X141 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X142 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X143 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X145 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X146 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X147 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X148 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X149 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X150 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X151 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X152 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X153 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X154 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X155 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X156 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X157 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X158 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X159 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X160 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X161 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X162 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X163 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X164 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X165 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X166 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X167 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X168 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X169 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X170 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X171 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X172 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X173 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X174 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X175 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X176 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X177 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X178 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X179 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X180 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X181 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X182 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X183 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X184 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X185 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X186 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X187 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X188 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X189 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X190 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X191 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X192 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X193 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X194 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X195 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X196 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X197 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X198 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X199 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X200 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X201 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X202 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X203 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X204 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X205 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X206 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X207 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X208 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X209 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X210 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X211 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X212 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X213 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X214 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X215 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X216 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X217 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X218 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X219 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X220 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X221 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X222 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X223 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X224 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X225 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X226 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X227 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X228 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X229 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X230 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X231 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X232 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X233 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X234 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X235 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X236 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X237 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X238 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X239 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X240 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X241 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X242 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X243 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X244 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X245 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X246 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X247 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X248 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X249 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X250 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X251 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X252 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X253 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X254 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X255 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X256 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X257 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X258 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X259 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X261 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X262 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X263 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X264 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X265 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X266 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X267 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X268 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X269 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X273 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X274 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X275 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X276 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X277 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X279 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X280 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X281 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X283 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X284 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X285 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X286 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X287 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X288 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X289 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X290 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X291 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X292 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X293 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X294 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X295 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X296 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X297 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X298 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X299 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X300 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X301 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X302 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X303 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X304 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X305 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X306 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X307 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X308 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X309 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X310 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X311 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X312 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X313 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X314 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X315 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X316 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X317 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X318 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X319 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X320 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X321 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X322 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X323 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X324 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X325 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X326 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X327 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X328 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X329 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X330 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X331 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X332 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X333 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X334 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X335 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X336 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X337 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X338 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X339 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X340 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X341 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X342 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X343 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X344 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X345 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X346 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X347 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X348 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X349 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X350 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X351 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X352 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X353 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X354 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X355 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X356 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X357 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X358 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X359 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X360 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X361 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X362 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X363 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X364 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X365 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X366 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X367 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X368 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X369 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X370 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X371 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X372 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X373 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X374 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X375 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X376 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X377 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X378 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X379 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X380 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X381 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X382 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X383 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X384 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X385 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X386 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X387 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X388 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X389 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X390 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X391 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X392 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X393 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X394 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X395 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X396 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X397 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X398 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X399 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X400 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X401 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X402 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X403 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X404 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X405 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X406 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X407 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X408 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X409 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X410 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X411 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X412 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X413 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X414 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X415 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X416 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X417 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X418 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X419 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X420 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X421 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X422 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X423 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X424 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X425 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X426 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X427 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X428 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X429 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X430 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X431 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X432 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X433 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X434 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X435 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X436 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X437 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X438 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X439 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X440 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X441 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X442 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X443 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X444 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X445 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X446 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X447 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X448 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X449 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X450 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X451 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X452 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X453 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X454 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X455 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X456 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X457 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X458 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X459 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X460 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X461 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X462 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X463 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X464 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X465 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X466 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X467 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X468 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X469 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X470 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X471 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X472 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X473 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X474 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X475 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X476 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X477 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X478 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X479 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X480 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X481 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X482 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X483 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X484 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X485 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X486 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X487 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X488 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X489 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X490 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X491 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X492 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X493 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X494 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X495 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X496 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X497 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X498 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X499 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X500 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X501 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X502 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X503 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X504 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X505 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X506 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X507 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X508 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X509 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X510 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X511 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X512 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X513 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X514 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X515 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X516 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X517 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X519 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X520 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X521 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X522 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X523 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X524 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X525 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X526 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X527 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X528 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X529 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X530 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X531 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X532 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X533 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X534 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X535 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X536 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X537 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X538 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X540 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X541 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X542 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X543 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X544 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X545 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X546 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X547 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X548 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X549 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X550 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X551 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X552 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X553 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X554 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X555 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X556 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X557 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X558 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X559 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X560 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X561 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X562 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X563 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X564 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X565 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X566 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X567 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X568 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X569 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X570 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X571 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X572 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X573 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X574 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X575 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X576 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X577 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X578 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X579 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X580 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X581 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X582 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X583 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X584 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X585 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X586 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X587 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X588 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X589 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X590 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X591 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X592 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X593 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X594 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X595 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X596 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X597 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X598 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X599 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X600 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X601 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X602 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X603 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X604 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X605 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X606 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X607 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X608 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X609 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X610 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X611 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X612 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X613 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X614 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X615 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X616 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X617 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X618 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X619 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X620 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X621 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X622 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X623 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X624 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X625 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X626 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X627 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X628 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X629 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X630 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X631 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X632 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X633 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X634 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X635 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X636 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X637 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X638 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X639 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X640 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X641 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X642 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X643 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X644 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X645 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X646 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X647 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X648 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X649 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X650 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X651 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X652 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X653 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X654 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X655 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X656 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X657 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X658 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X659 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X660 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X661 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X662 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X663 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X664 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X665 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X666 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X667 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X668 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X669 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X670 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X671 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X672 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X673 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X674 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X675 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X676 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X677 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X678 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X679 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X680 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X681 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X682 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X683 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X684 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X685 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X686 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X687 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X688 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X689 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X690 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X691 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X692 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X693 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X694 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X695 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X696 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X697 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X698 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X699 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X700 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X701 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X702 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X703 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X704 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X705 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X706 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X707 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X708 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X709 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X710 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X711 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X712 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X713 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X714 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X715 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X716 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X717 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X718 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X719 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X720 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X721 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X722 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X723 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X724 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X725 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X726 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X727 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X728 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X729 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X730 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X731 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X732 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X733 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X734 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X735 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X736 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X737 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X738 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X739 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X740 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X741 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X742 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X743 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X744 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X745 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X746 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X747 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X748 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X749 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X750 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X751 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X752 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X753 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X754 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X755 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X756 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X757 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X758 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X759 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X760 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X761 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X762 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X763 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X764 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X765 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X766 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X767 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X768 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X769 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X770 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X771 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X772 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X773 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X774 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X775 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X776 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X777 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X778 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X779 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X780 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X781 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X782 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X783 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X784 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X785 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X786 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X787 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X788 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X789 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X790 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X791 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X792 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X793 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X794 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X795 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X796 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X797 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X798 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X799 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X800 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X801 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X802 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X803 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X804 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X805 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X806 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X807 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X808 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X809 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X810 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X811 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X812 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X813 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X814 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X815 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X816 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X817 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X818 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X819 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X820 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X821 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X822 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X823 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X824 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X825 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X826 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X827 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X828 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X829 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X830 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X831 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X832 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X833 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X834 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X835 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X836 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X837 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X838 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X839 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X840 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X841 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X842 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X843 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X844 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X845 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X846 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X847 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X848 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X849 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X850 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X851 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X852 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X853 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X854 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X855 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X856 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X857 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X858 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X859 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X860 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X861 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X862 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X863 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X864 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X865 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X866 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X867 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X868 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X869 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X870 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X871 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X872 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X873 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X874 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X875 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X876 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X877 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X878 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X879 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X880 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X881 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X882 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X883 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X884 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X885 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X886 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X887 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X888 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X889 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X890 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X891 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X892 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X893 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X894 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X895 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X896 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X897 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X898 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X899 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X900 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X901 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X902 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X903 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X904 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X905 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X906 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X907 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X908 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X909 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X910 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X911 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X912 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X913 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X914 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X915 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X916 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X917 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X918 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X919 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X920 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X921 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X922 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X923 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X924 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X925 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X926 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X927 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X928 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X929 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X930 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X931 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X932 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X933 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X934 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X935 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X936 cmirror_out m1_250_8900# m1_370_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X937 m1_370_11400# m1_250_8900# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X938 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X939 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X940 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X941 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X942 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X943 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X944 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X945 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X946 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X947 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X948 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X949 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X950 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X951 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X952 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X953 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X954 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X955 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X956 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X957 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X958 cmirror_out m1_1850_8370# m1_2350_11400# cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X959 m1_2350_11400# m1_1850_8370# cmirror_out cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X960 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X961 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X962 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X963 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X964 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X965 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X966 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X967 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X968 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X969 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X970 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X971 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X972 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X973 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X974 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X975 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X976 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X977 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X978 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X979 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X980 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X981 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X982 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X983 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X984 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X985 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X986 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X987 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X988 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X989 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X990 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X991 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X992 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X993 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X994 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X995 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X996 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X997 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X998 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X999 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1000 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1001 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1002 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1003 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1004 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1005 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1006 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1007 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1008 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1009 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1010 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1011 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1012 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1013 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1014 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1015 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1016 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1017 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1018 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1019 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1020 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1021 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1022 cmirror_out outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1023 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1024 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1025 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1026 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1027 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1028 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1029 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1030 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1031 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1032 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1033 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1034 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1035 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1036 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1037 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1038 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1039 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1040 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1041 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1042 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1043 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1044 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1045 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1046 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1047 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1048 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1049 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1050 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1051 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1052 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1053 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1054 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1055 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1056 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1057 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1058 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1059 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1060 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1061 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1062 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1063 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1064 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1065 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1066 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1067 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1068 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1069 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1070 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1071 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1072 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1073 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1074 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1075 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1076 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1077 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1078 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1079 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1080 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1081 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1082 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1083 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1084 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1085 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1086 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1087 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1088 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1089 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1090 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1091 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1092 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1093 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1094 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1095 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1096 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1097 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1098 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1099 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1100 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1101 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1102 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1103 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1104 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1105 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1106 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1107 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1108 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1109 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1110 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1111 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1112 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1113 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1114 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1115 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1116 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1117 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1118 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1119 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1120 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1121 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1122 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1123 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1124 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1125 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1126 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1127 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1128 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1129 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1130 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1131 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1132 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1133 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1134 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1135 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1136 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1137 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1138 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1139 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1140 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1141 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1142 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1143 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1144 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1145 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1146 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1147 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1148 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1149 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1150 VN outd_cmirror_64t_4/m1_0_80# m2_7240_7300# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1151 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
