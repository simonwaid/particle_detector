* SPICE3 file created from esd-array.ext - technology: sky130A

D0 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D1 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D2 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D3 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D4 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D5 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D6 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D7 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D8 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D9 m1_n9140_490# w_n2010_1280# sky130_fd_pr__diode_pd2nw_11v0 pj=8e+06u area=4e+12p
D10 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D11 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D12 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D13 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D14 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D15 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D16 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D17 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D18 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
D19 VSUBS m1_n9140_490# sky130_fd_pr__diode_pw2nd_11v0 pj=8e+06u area=4e+12p
