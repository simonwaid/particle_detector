magic
tech sky130A
magscale 1 2
timestamp 1645462850
<< pwell >>
rect -6457 -1119 6457 1119
<< nmos >>
rect -6261 109 -5061 909
rect -5003 109 -3803 909
rect -3745 109 -2545 909
rect -2487 109 -1287 909
rect -1229 109 -29 909
rect 29 109 1229 909
rect 1287 109 2487 909
rect 2545 109 3745 909
rect 3803 109 5003 909
rect 5061 109 6261 909
rect -6261 -909 -5061 -109
rect -5003 -909 -3803 -109
rect -3745 -909 -2545 -109
rect -2487 -909 -1287 -109
rect -1229 -909 -29 -109
rect 29 -909 1229 -109
rect 1287 -909 2487 -109
rect 2545 -909 3745 -109
rect 3803 -909 5003 -109
rect 5061 -909 6261 -109
<< ndiff >>
rect -6319 897 -6261 909
rect -6319 121 -6307 897
rect -6273 121 -6261 897
rect -6319 109 -6261 121
rect -5061 897 -5003 909
rect -5061 121 -5049 897
rect -5015 121 -5003 897
rect -5061 109 -5003 121
rect -3803 897 -3745 909
rect -3803 121 -3791 897
rect -3757 121 -3745 897
rect -3803 109 -3745 121
rect -2545 897 -2487 909
rect -2545 121 -2533 897
rect -2499 121 -2487 897
rect -2545 109 -2487 121
rect -1287 897 -1229 909
rect -1287 121 -1275 897
rect -1241 121 -1229 897
rect -1287 109 -1229 121
rect -29 897 29 909
rect -29 121 -17 897
rect 17 121 29 897
rect -29 109 29 121
rect 1229 897 1287 909
rect 1229 121 1241 897
rect 1275 121 1287 897
rect 1229 109 1287 121
rect 2487 897 2545 909
rect 2487 121 2499 897
rect 2533 121 2545 897
rect 2487 109 2545 121
rect 3745 897 3803 909
rect 3745 121 3757 897
rect 3791 121 3803 897
rect 3745 109 3803 121
rect 5003 897 5061 909
rect 5003 121 5015 897
rect 5049 121 5061 897
rect 5003 109 5061 121
rect 6261 897 6319 909
rect 6261 121 6273 897
rect 6307 121 6319 897
rect 6261 109 6319 121
rect -6319 -121 -6261 -109
rect -6319 -897 -6307 -121
rect -6273 -897 -6261 -121
rect -6319 -909 -6261 -897
rect -5061 -121 -5003 -109
rect -5061 -897 -5049 -121
rect -5015 -897 -5003 -121
rect -5061 -909 -5003 -897
rect -3803 -121 -3745 -109
rect -3803 -897 -3791 -121
rect -3757 -897 -3745 -121
rect -3803 -909 -3745 -897
rect -2545 -121 -2487 -109
rect -2545 -897 -2533 -121
rect -2499 -897 -2487 -121
rect -2545 -909 -2487 -897
rect -1287 -121 -1229 -109
rect -1287 -897 -1275 -121
rect -1241 -897 -1229 -121
rect -1287 -909 -1229 -897
rect -29 -121 29 -109
rect -29 -897 -17 -121
rect 17 -897 29 -121
rect -29 -909 29 -897
rect 1229 -121 1287 -109
rect 1229 -897 1241 -121
rect 1275 -897 1287 -121
rect 1229 -909 1287 -897
rect 2487 -121 2545 -109
rect 2487 -897 2499 -121
rect 2533 -897 2545 -121
rect 2487 -909 2545 -897
rect 3745 -121 3803 -109
rect 3745 -897 3757 -121
rect 3791 -897 3803 -121
rect 3745 -909 3803 -897
rect 5003 -121 5061 -109
rect 5003 -897 5015 -121
rect 5049 -897 5061 -121
rect 5003 -909 5061 -897
rect 6261 -121 6319 -109
rect 6261 -897 6273 -121
rect 6307 -897 6319 -121
rect 6261 -909 6319 -897
<< ndiffc >>
rect -6307 121 -6273 897
rect -5049 121 -5015 897
rect -3791 121 -3757 897
rect -2533 121 -2499 897
rect -1275 121 -1241 897
rect -17 121 17 897
rect 1241 121 1275 897
rect 2499 121 2533 897
rect 3757 121 3791 897
rect 5015 121 5049 897
rect 6273 121 6307 897
rect -6307 -897 -6273 -121
rect -5049 -897 -5015 -121
rect -3791 -897 -3757 -121
rect -2533 -897 -2499 -121
rect -1275 -897 -1241 -121
rect -17 -897 17 -121
rect 1241 -897 1275 -121
rect 2499 -897 2533 -121
rect 3757 -897 3791 -121
rect 5015 -897 5049 -121
rect 6273 -897 6307 -121
<< psubdiff >>
rect -6421 1049 -6325 1083
rect 6325 1049 6421 1083
rect -6421 987 -6387 1049
rect 6387 987 6421 1049
rect -6421 -1049 -6387 -987
rect 6387 -1049 6421 -987
rect -6421 -1083 -6325 -1049
rect 6325 -1083 6421 -1049
<< psubdiffcont >>
rect -6325 1049 6325 1083
rect -6421 -987 -6387 987
rect 6387 -987 6421 987
rect -6325 -1083 6325 -1049
<< poly >>
rect -6261 981 -5061 997
rect -6261 947 -6245 981
rect -5077 947 -5061 981
rect -6261 909 -5061 947
rect -5003 981 -3803 997
rect -5003 947 -4987 981
rect -3819 947 -3803 981
rect -5003 909 -3803 947
rect -3745 981 -2545 997
rect -3745 947 -3729 981
rect -2561 947 -2545 981
rect -3745 909 -2545 947
rect -2487 981 -1287 997
rect -2487 947 -2471 981
rect -1303 947 -1287 981
rect -2487 909 -1287 947
rect -1229 981 -29 997
rect -1229 947 -1213 981
rect -45 947 -29 981
rect -1229 909 -29 947
rect 29 981 1229 997
rect 29 947 45 981
rect 1213 947 1229 981
rect 29 909 1229 947
rect 1287 981 2487 997
rect 1287 947 1303 981
rect 2471 947 2487 981
rect 1287 909 2487 947
rect 2545 981 3745 997
rect 2545 947 2561 981
rect 3729 947 3745 981
rect 2545 909 3745 947
rect 3803 981 5003 997
rect 3803 947 3819 981
rect 4987 947 5003 981
rect 3803 909 5003 947
rect 5061 981 6261 997
rect 5061 947 5077 981
rect 6245 947 6261 981
rect 5061 909 6261 947
rect -6261 71 -5061 109
rect -6261 37 -6245 71
rect -5077 37 -5061 71
rect -6261 21 -5061 37
rect -5003 71 -3803 109
rect -5003 37 -4987 71
rect -3819 37 -3803 71
rect -5003 21 -3803 37
rect -3745 71 -2545 109
rect -3745 37 -3729 71
rect -2561 37 -2545 71
rect -3745 21 -2545 37
rect -2487 71 -1287 109
rect -2487 37 -2471 71
rect -1303 37 -1287 71
rect -2487 21 -1287 37
rect -1229 71 -29 109
rect -1229 37 -1213 71
rect -45 37 -29 71
rect -1229 21 -29 37
rect 29 71 1229 109
rect 29 37 45 71
rect 1213 37 1229 71
rect 29 21 1229 37
rect 1287 71 2487 109
rect 1287 37 1303 71
rect 2471 37 2487 71
rect 1287 21 2487 37
rect 2545 71 3745 109
rect 2545 37 2561 71
rect 3729 37 3745 71
rect 2545 21 3745 37
rect 3803 71 5003 109
rect 3803 37 3819 71
rect 4987 37 5003 71
rect 3803 21 5003 37
rect 5061 71 6261 109
rect 5061 37 5077 71
rect 6245 37 6261 71
rect 5061 21 6261 37
rect -6261 -37 -5061 -21
rect -6261 -71 -6245 -37
rect -5077 -71 -5061 -37
rect -6261 -109 -5061 -71
rect -5003 -37 -3803 -21
rect -5003 -71 -4987 -37
rect -3819 -71 -3803 -37
rect -5003 -109 -3803 -71
rect -3745 -37 -2545 -21
rect -3745 -71 -3729 -37
rect -2561 -71 -2545 -37
rect -3745 -109 -2545 -71
rect -2487 -37 -1287 -21
rect -2487 -71 -2471 -37
rect -1303 -71 -1287 -37
rect -2487 -109 -1287 -71
rect -1229 -37 -29 -21
rect -1229 -71 -1213 -37
rect -45 -71 -29 -37
rect -1229 -109 -29 -71
rect 29 -37 1229 -21
rect 29 -71 45 -37
rect 1213 -71 1229 -37
rect 29 -109 1229 -71
rect 1287 -37 2487 -21
rect 1287 -71 1303 -37
rect 2471 -71 2487 -37
rect 1287 -109 2487 -71
rect 2545 -37 3745 -21
rect 2545 -71 2561 -37
rect 3729 -71 3745 -37
rect 2545 -109 3745 -71
rect 3803 -37 5003 -21
rect 3803 -71 3819 -37
rect 4987 -71 5003 -37
rect 3803 -109 5003 -71
rect 5061 -37 6261 -21
rect 5061 -71 5077 -37
rect 6245 -71 6261 -37
rect 5061 -109 6261 -71
rect -6261 -947 -5061 -909
rect -6261 -981 -6245 -947
rect -5077 -981 -5061 -947
rect -6261 -997 -5061 -981
rect -5003 -947 -3803 -909
rect -5003 -981 -4987 -947
rect -3819 -981 -3803 -947
rect -5003 -997 -3803 -981
rect -3745 -947 -2545 -909
rect -3745 -981 -3729 -947
rect -2561 -981 -2545 -947
rect -3745 -997 -2545 -981
rect -2487 -947 -1287 -909
rect -2487 -981 -2471 -947
rect -1303 -981 -1287 -947
rect -2487 -997 -1287 -981
rect -1229 -947 -29 -909
rect -1229 -981 -1213 -947
rect -45 -981 -29 -947
rect -1229 -997 -29 -981
rect 29 -947 1229 -909
rect 29 -981 45 -947
rect 1213 -981 1229 -947
rect 29 -997 1229 -981
rect 1287 -947 2487 -909
rect 1287 -981 1303 -947
rect 2471 -981 2487 -947
rect 1287 -997 2487 -981
rect 2545 -947 3745 -909
rect 2545 -981 2561 -947
rect 3729 -981 3745 -947
rect 2545 -997 3745 -981
rect 3803 -947 5003 -909
rect 3803 -981 3819 -947
rect 4987 -981 5003 -947
rect 3803 -997 5003 -981
rect 5061 -947 6261 -909
rect 5061 -981 5077 -947
rect 6245 -981 6261 -947
rect 5061 -997 6261 -981
<< polycont >>
rect -6245 947 -5077 981
rect -4987 947 -3819 981
rect -3729 947 -2561 981
rect -2471 947 -1303 981
rect -1213 947 -45 981
rect 45 947 1213 981
rect 1303 947 2471 981
rect 2561 947 3729 981
rect 3819 947 4987 981
rect 5077 947 6245 981
rect -6245 37 -5077 71
rect -4987 37 -3819 71
rect -3729 37 -2561 71
rect -2471 37 -1303 71
rect -1213 37 -45 71
rect 45 37 1213 71
rect 1303 37 2471 71
rect 2561 37 3729 71
rect 3819 37 4987 71
rect 5077 37 6245 71
rect -6245 -71 -5077 -37
rect -4987 -71 -3819 -37
rect -3729 -71 -2561 -37
rect -2471 -71 -1303 -37
rect -1213 -71 -45 -37
rect 45 -71 1213 -37
rect 1303 -71 2471 -37
rect 2561 -71 3729 -37
rect 3819 -71 4987 -37
rect 5077 -71 6245 -37
rect -6245 -981 -5077 -947
rect -4987 -981 -3819 -947
rect -3729 -981 -2561 -947
rect -2471 -981 -1303 -947
rect -1213 -981 -45 -947
rect 45 -981 1213 -947
rect 1303 -981 2471 -947
rect 2561 -981 3729 -947
rect 3819 -981 4987 -947
rect 5077 -981 6245 -947
<< locali >>
rect -6421 1049 -6325 1083
rect 6325 1049 6421 1083
rect -6421 987 -6387 1049
rect 6387 987 6421 1049
rect -6261 947 -6245 981
rect -5077 947 -5061 981
rect -5003 947 -4987 981
rect -3819 947 -3803 981
rect -3745 947 -3729 981
rect -2561 947 -2545 981
rect -2487 947 -2471 981
rect -1303 947 -1287 981
rect -1229 947 -1213 981
rect -45 947 -29 981
rect 29 947 45 981
rect 1213 947 1229 981
rect 1287 947 1303 981
rect 2471 947 2487 981
rect 2545 947 2561 981
rect 3729 947 3745 981
rect 3803 947 3819 981
rect 4987 947 5003 981
rect 5061 947 5077 981
rect 6245 947 6261 981
rect -6307 897 -6273 913
rect -6307 105 -6273 121
rect -5049 897 -5015 913
rect -5049 105 -5015 121
rect -3791 897 -3757 913
rect -3791 105 -3757 121
rect -2533 897 -2499 913
rect -2533 105 -2499 121
rect -1275 897 -1241 913
rect -1275 105 -1241 121
rect -17 897 17 913
rect -17 105 17 121
rect 1241 897 1275 913
rect 1241 105 1275 121
rect 2499 897 2533 913
rect 2499 105 2533 121
rect 3757 897 3791 913
rect 3757 105 3791 121
rect 5015 897 5049 913
rect 5015 105 5049 121
rect 6273 897 6307 913
rect 6273 105 6307 121
rect -6261 37 -6245 71
rect -5077 37 -5061 71
rect -5003 37 -4987 71
rect -3819 37 -3803 71
rect -3745 37 -3729 71
rect -2561 37 -2545 71
rect -2487 37 -2471 71
rect -1303 37 -1287 71
rect -1229 37 -1213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1213 37 1229 71
rect 1287 37 1303 71
rect 2471 37 2487 71
rect 2545 37 2561 71
rect 3729 37 3745 71
rect 3803 37 3819 71
rect 4987 37 5003 71
rect 5061 37 5077 71
rect 6245 37 6261 71
rect -6261 -71 -6245 -37
rect -5077 -71 -5061 -37
rect -5003 -71 -4987 -37
rect -3819 -71 -3803 -37
rect -3745 -71 -3729 -37
rect -2561 -71 -2545 -37
rect -2487 -71 -2471 -37
rect -1303 -71 -1287 -37
rect -1229 -71 -1213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1213 -71 1229 -37
rect 1287 -71 1303 -37
rect 2471 -71 2487 -37
rect 2545 -71 2561 -37
rect 3729 -71 3745 -37
rect 3803 -71 3819 -37
rect 4987 -71 5003 -37
rect 5061 -71 5077 -37
rect 6245 -71 6261 -37
rect -6307 -121 -6273 -105
rect -6307 -913 -6273 -897
rect -5049 -121 -5015 -105
rect -5049 -913 -5015 -897
rect -3791 -121 -3757 -105
rect -3791 -913 -3757 -897
rect -2533 -121 -2499 -105
rect -2533 -913 -2499 -897
rect -1275 -121 -1241 -105
rect -1275 -913 -1241 -897
rect -17 -121 17 -105
rect -17 -913 17 -897
rect 1241 -121 1275 -105
rect 1241 -913 1275 -897
rect 2499 -121 2533 -105
rect 2499 -913 2533 -897
rect 3757 -121 3791 -105
rect 3757 -913 3791 -897
rect 5015 -121 5049 -105
rect 5015 -913 5049 -897
rect 6273 -121 6307 -105
rect 6273 -913 6307 -897
rect -6261 -981 -6245 -947
rect -5077 -981 -5061 -947
rect -5003 -981 -4987 -947
rect -3819 -981 -3803 -947
rect -3745 -981 -3729 -947
rect -2561 -981 -2545 -947
rect -2487 -981 -2471 -947
rect -1303 -981 -1287 -947
rect -1229 -981 -1213 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 1213 -981 1229 -947
rect 1287 -981 1303 -947
rect 2471 -981 2487 -947
rect 2545 -981 2561 -947
rect 3729 -981 3745 -947
rect 3803 -981 3819 -947
rect 4987 -981 5003 -947
rect 5061 -981 5077 -947
rect 6245 -981 6261 -947
rect -6421 -1049 -6387 -987
rect 6387 -1049 6421 -987
rect -6421 -1083 -6325 -1049
rect 6325 -1083 6421 -1049
<< viali >>
rect -6245 947 -5077 981
rect -4987 947 -3819 981
rect -3729 947 -2561 981
rect -2471 947 -1303 981
rect -1213 947 -45 981
rect 45 947 1213 981
rect 1303 947 2471 981
rect 2561 947 3729 981
rect 3819 947 4987 981
rect 5077 947 6245 981
rect -6307 121 -6273 897
rect -5049 121 -5015 897
rect -3791 121 -3757 897
rect -2533 121 -2499 897
rect -1275 121 -1241 897
rect -17 121 17 897
rect 1241 121 1275 897
rect 2499 121 2533 897
rect 3757 121 3791 897
rect 5015 121 5049 897
rect 6273 121 6307 897
rect -6245 37 -5077 71
rect -4987 37 -3819 71
rect -3729 37 -2561 71
rect -2471 37 -1303 71
rect -1213 37 -45 71
rect 45 37 1213 71
rect 1303 37 2471 71
rect 2561 37 3729 71
rect 3819 37 4987 71
rect 5077 37 6245 71
rect -6245 -71 -5077 -37
rect -4987 -71 -3819 -37
rect -3729 -71 -2561 -37
rect -2471 -71 -1303 -37
rect -1213 -71 -45 -37
rect 45 -71 1213 -37
rect 1303 -71 2471 -37
rect 2561 -71 3729 -37
rect 3819 -71 4987 -37
rect 5077 -71 6245 -37
rect -6307 -897 -6273 -121
rect -5049 -897 -5015 -121
rect -3791 -897 -3757 -121
rect -2533 -897 -2499 -121
rect -1275 -897 -1241 -121
rect -17 -897 17 -121
rect 1241 -897 1275 -121
rect 2499 -897 2533 -121
rect 3757 -897 3791 -121
rect 5015 -897 5049 -121
rect 6273 -897 6307 -121
rect -6245 -981 -5077 -947
rect -4987 -981 -3819 -947
rect -3729 -981 -2561 -947
rect -2471 -981 -1303 -947
rect -1213 -981 -45 -947
rect 45 -981 1213 -947
rect 1303 -981 2471 -947
rect 2561 -981 3729 -947
rect 3819 -981 4987 -947
rect 5077 -981 6245 -947
<< metal1 >>
rect -6257 981 -5065 987
rect -6257 947 -6245 981
rect -5077 947 -5065 981
rect -6257 941 -5065 947
rect -4999 981 -3807 987
rect -4999 947 -4987 981
rect -3819 947 -3807 981
rect -4999 941 -3807 947
rect -3741 981 -2549 987
rect -3741 947 -3729 981
rect -2561 947 -2549 981
rect -3741 941 -2549 947
rect -2483 981 -1291 987
rect -2483 947 -2471 981
rect -1303 947 -1291 981
rect -2483 941 -1291 947
rect -1225 981 -33 987
rect -1225 947 -1213 981
rect -45 947 -33 981
rect -1225 941 -33 947
rect 33 981 1225 987
rect 33 947 45 981
rect 1213 947 1225 981
rect 33 941 1225 947
rect 1291 981 2483 987
rect 1291 947 1303 981
rect 2471 947 2483 981
rect 1291 941 2483 947
rect 2549 981 3741 987
rect 2549 947 2561 981
rect 3729 947 3741 981
rect 2549 941 3741 947
rect 3807 981 4999 987
rect 3807 947 3819 981
rect 4987 947 4999 981
rect 3807 941 4999 947
rect 5065 981 6257 987
rect 5065 947 5077 981
rect 6245 947 6257 981
rect 5065 941 6257 947
rect -6313 897 -6267 909
rect -6313 121 -6307 897
rect -6273 121 -6267 897
rect -6313 109 -6267 121
rect -5055 897 -5009 909
rect -5055 121 -5049 897
rect -5015 121 -5009 897
rect -5055 109 -5009 121
rect -3797 897 -3751 909
rect -3797 121 -3791 897
rect -3757 121 -3751 897
rect -3797 109 -3751 121
rect -2539 897 -2493 909
rect -2539 121 -2533 897
rect -2499 121 -2493 897
rect -2539 109 -2493 121
rect -1281 897 -1235 909
rect -1281 121 -1275 897
rect -1241 121 -1235 897
rect -1281 109 -1235 121
rect -23 897 23 909
rect -23 121 -17 897
rect 17 121 23 897
rect -23 109 23 121
rect 1235 897 1281 909
rect 1235 121 1241 897
rect 1275 121 1281 897
rect 1235 109 1281 121
rect 2493 897 2539 909
rect 2493 121 2499 897
rect 2533 121 2539 897
rect 2493 109 2539 121
rect 3751 897 3797 909
rect 3751 121 3757 897
rect 3791 121 3797 897
rect 3751 109 3797 121
rect 5009 897 5055 909
rect 5009 121 5015 897
rect 5049 121 5055 897
rect 5009 109 5055 121
rect 6267 897 6313 909
rect 6267 121 6273 897
rect 6307 121 6313 897
rect 6267 109 6313 121
rect -6257 71 -5065 77
rect -6257 37 -6245 71
rect -5077 37 -5065 71
rect -6257 31 -5065 37
rect -4999 71 -3807 77
rect -4999 37 -4987 71
rect -3819 37 -3807 71
rect -4999 31 -3807 37
rect -3741 71 -2549 77
rect -3741 37 -3729 71
rect -2561 37 -2549 71
rect -3741 31 -2549 37
rect -2483 71 -1291 77
rect -2483 37 -2471 71
rect -1303 37 -1291 71
rect -2483 31 -1291 37
rect -1225 71 -33 77
rect -1225 37 -1213 71
rect -45 37 -33 71
rect -1225 31 -33 37
rect 33 71 1225 77
rect 33 37 45 71
rect 1213 37 1225 71
rect 33 31 1225 37
rect 1291 71 2483 77
rect 1291 37 1303 71
rect 2471 37 2483 71
rect 1291 31 2483 37
rect 2549 71 3741 77
rect 2549 37 2561 71
rect 3729 37 3741 71
rect 2549 31 3741 37
rect 3807 71 4999 77
rect 3807 37 3819 71
rect 4987 37 4999 71
rect 3807 31 4999 37
rect 5065 71 6257 77
rect 5065 37 5077 71
rect 6245 37 6257 71
rect 5065 31 6257 37
rect -6257 -37 -5065 -31
rect -6257 -71 -6245 -37
rect -5077 -71 -5065 -37
rect -6257 -77 -5065 -71
rect -4999 -37 -3807 -31
rect -4999 -71 -4987 -37
rect -3819 -71 -3807 -37
rect -4999 -77 -3807 -71
rect -3741 -37 -2549 -31
rect -3741 -71 -3729 -37
rect -2561 -71 -2549 -37
rect -3741 -77 -2549 -71
rect -2483 -37 -1291 -31
rect -2483 -71 -2471 -37
rect -1303 -71 -1291 -37
rect -2483 -77 -1291 -71
rect -1225 -37 -33 -31
rect -1225 -71 -1213 -37
rect -45 -71 -33 -37
rect -1225 -77 -33 -71
rect 33 -37 1225 -31
rect 33 -71 45 -37
rect 1213 -71 1225 -37
rect 33 -77 1225 -71
rect 1291 -37 2483 -31
rect 1291 -71 1303 -37
rect 2471 -71 2483 -37
rect 1291 -77 2483 -71
rect 2549 -37 3741 -31
rect 2549 -71 2561 -37
rect 3729 -71 3741 -37
rect 2549 -77 3741 -71
rect 3807 -37 4999 -31
rect 3807 -71 3819 -37
rect 4987 -71 4999 -37
rect 3807 -77 4999 -71
rect 5065 -37 6257 -31
rect 5065 -71 5077 -37
rect 6245 -71 6257 -37
rect 5065 -77 6257 -71
rect -6313 -121 -6267 -109
rect -6313 -897 -6307 -121
rect -6273 -897 -6267 -121
rect -6313 -909 -6267 -897
rect -5055 -121 -5009 -109
rect -5055 -897 -5049 -121
rect -5015 -897 -5009 -121
rect -5055 -909 -5009 -897
rect -3797 -121 -3751 -109
rect -3797 -897 -3791 -121
rect -3757 -897 -3751 -121
rect -3797 -909 -3751 -897
rect -2539 -121 -2493 -109
rect -2539 -897 -2533 -121
rect -2499 -897 -2493 -121
rect -2539 -909 -2493 -897
rect -1281 -121 -1235 -109
rect -1281 -897 -1275 -121
rect -1241 -897 -1235 -121
rect -1281 -909 -1235 -897
rect -23 -121 23 -109
rect -23 -897 -17 -121
rect 17 -897 23 -121
rect -23 -909 23 -897
rect 1235 -121 1281 -109
rect 1235 -897 1241 -121
rect 1275 -897 1281 -121
rect 1235 -909 1281 -897
rect 2493 -121 2539 -109
rect 2493 -897 2499 -121
rect 2533 -897 2539 -121
rect 2493 -909 2539 -897
rect 3751 -121 3797 -109
rect 3751 -897 3757 -121
rect 3791 -897 3797 -121
rect 3751 -909 3797 -897
rect 5009 -121 5055 -109
rect 5009 -897 5015 -121
rect 5049 -897 5055 -121
rect 5009 -909 5055 -897
rect 6267 -121 6313 -109
rect 6267 -897 6273 -121
rect 6307 -897 6313 -121
rect 6267 -909 6313 -897
rect -6257 -947 -5065 -941
rect -6257 -981 -6245 -947
rect -5077 -981 -5065 -947
rect -6257 -987 -5065 -981
rect -4999 -947 -3807 -941
rect -4999 -981 -4987 -947
rect -3819 -981 -3807 -947
rect -4999 -987 -3807 -981
rect -3741 -947 -2549 -941
rect -3741 -981 -3729 -947
rect -2561 -981 -2549 -947
rect -3741 -987 -2549 -981
rect -2483 -947 -1291 -941
rect -2483 -981 -2471 -947
rect -1303 -981 -1291 -947
rect -2483 -987 -1291 -981
rect -1225 -947 -33 -941
rect -1225 -981 -1213 -947
rect -45 -981 -33 -947
rect -1225 -987 -33 -981
rect 33 -947 1225 -941
rect 33 -981 45 -947
rect 1213 -981 1225 -947
rect 33 -987 1225 -981
rect 1291 -947 2483 -941
rect 1291 -981 1303 -947
rect 2471 -981 2483 -947
rect 1291 -987 2483 -981
rect 2549 -947 3741 -941
rect 2549 -981 2561 -947
rect 3729 -981 3741 -947
rect 2549 -987 3741 -981
rect 3807 -947 4999 -941
rect 3807 -981 3819 -947
rect 4987 -981 4999 -947
rect 3807 -987 4999 -981
rect 5065 -947 6257 -941
rect 5065 -981 5077 -947
rect 6245 -981 6257 -947
rect 5065 -987 6257 -981
<< properties >>
string FIXED_BBOX -6404 -1066 6404 1066
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 6 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
