magic
tech sky130A
magscale 1 2
timestamp 1646400034
<< nwell >>
rect -1083 -755 1083 755
<< pmos >>
rect -887 336 -487 536
rect -429 336 -29 536
rect 29 336 429 536
rect 487 336 887 536
rect -887 -100 -487 100
rect -429 -100 -29 100
rect 29 -100 429 100
rect 487 -100 887 100
rect -887 -536 -487 -336
rect -429 -536 -29 -336
rect 29 -536 429 -336
rect 487 -536 887 -336
<< pdiff >>
rect -945 524 -887 536
rect -945 348 -933 524
rect -899 348 -887 524
rect -945 336 -887 348
rect -487 524 -429 536
rect -487 348 -475 524
rect -441 348 -429 524
rect -487 336 -429 348
rect -29 524 29 536
rect -29 348 -17 524
rect 17 348 29 524
rect -29 336 29 348
rect 429 524 487 536
rect 429 348 441 524
rect 475 348 487 524
rect 429 336 487 348
rect 887 524 945 536
rect 887 348 899 524
rect 933 348 945 524
rect 887 336 945 348
rect -945 88 -887 100
rect -945 -88 -933 88
rect -899 -88 -887 88
rect -945 -100 -887 -88
rect -487 88 -429 100
rect -487 -88 -475 88
rect -441 -88 -429 88
rect -487 -100 -429 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 429 88 487 100
rect 429 -88 441 88
rect 475 -88 487 88
rect 429 -100 487 -88
rect 887 88 945 100
rect 887 -88 899 88
rect 933 -88 945 88
rect 887 -100 945 -88
rect -945 -348 -887 -336
rect -945 -524 -933 -348
rect -899 -524 -887 -348
rect -945 -536 -887 -524
rect -487 -348 -429 -336
rect -487 -524 -475 -348
rect -441 -524 -429 -348
rect -487 -536 -429 -524
rect -29 -348 29 -336
rect -29 -524 -17 -348
rect 17 -524 29 -348
rect -29 -536 29 -524
rect 429 -348 487 -336
rect 429 -524 441 -348
rect 475 -524 487 -348
rect 429 -536 487 -524
rect 887 -348 945 -336
rect 887 -524 899 -348
rect 933 -524 945 -348
rect 887 -536 945 -524
<< pdiffc >>
rect -933 348 -899 524
rect -475 348 -441 524
rect -17 348 17 524
rect 441 348 475 524
rect 899 348 933 524
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect -933 -524 -899 -348
rect -475 -524 -441 -348
rect -17 -524 17 -348
rect 441 -524 475 -348
rect 899 -524 933 -348
<< nsubdiff >>
rect -1047 685 -951 719
rect 951 685 1047 719
rect -1047 623 -1013 685
rect 1013 623 1047 685
rect -1047 -685 -1013 -623
rect 1013 -685 1047 -623
rect -1047 -719 -951 -685
rect 951 -719 1047 -685
<< nsubdiffcont >>
rect -951 685 951 719
rect -1047 -623 -1013 623
rect 1013 -623 1047 623
rect -951 -719 951 -685
<< poly >>
rect -887 617 -487 633
rect -887 583 -871 617
rect -503 583 -487 617
rect -887 536 -487 583
rect -429 617 -29 633
rect -429 583 -413 617
rect -45 583 -29 617
rect -429 536 -29 583
rect 29 617 429 633
rect 29 583 45 617
rect 413 583 429 617
rect 29 536 429 583
rect 487 617 887 633
rect 487 583 503 617
rect 871 583 887 617
rect 487 536 887 583
rect -887 289 -487 336
rect -887 255 -871 289
rect -503 255 -487 289
rect -887 239 -487 255
rect -429 289 -29 336
rect -429 255 -413 289
rect -45 255 -29 289
rect -429 239 -29 255
rect 29 289 429 336
rect 29 255 45 289
rect 413 255 429 289
rect 29 239 429 255
rect 487 289 887 336
rect 487 255 503 289
rect 871 255 887 289
rect 487 239 887 255
rect -887 181 -487 197
rect -887 147 -871 181
rect -503 147 -487 181
rect -887 100 -487 147
rect -429 181 -29 197
rect -429 147 -413 181
rect -45 147 -29 181
rect -429 100 -29 147
rect 29 181 429 197
rect 29 147 45 181
rect 413 147 429 181
rect 29 100 429 147
rect 487 181 887 197
rect 487 147 503 181
rect 871 147 887 181
rect 487 100 887 147
rect -887 -147 -487 -100
rect -887 -181 -871 -147
rect -503 -181 -487 -147
rect -887 -197 -487 -181
rect -429 -147 -29 -100
rect -429 -181 -413 -147
rect -45 -181 -29 -147
rect -429 -197 -29 -181
rect 29 -147 429 -100
rect 29 -181 45 -147
rect 413 -181 429 -147
rect 29 -197 429 -181
rect 487 -147 887 -100
rect 487 -181 503 -147
rect 871 -181 887 -147
rect 487 -197 887 -181
rect -887 -255 -487 -239
rect -887 -289 -871 -255
rect -503 -289 -487 -255
rect -887 -336 -487 -289
rect -429 -255 -29 -239
rect -429 -289 -413 -255
rect -45 -289 -29 -255
rect -429 -336 -29 -289
rect 29 -255 429 -239
rect 29 -289 45 -255
rect 413 -289 429 -255
rect 29 -336 429 -289
rect 487 -255 887 -239
rect 487 -289 503 -255
rect 871 -289 887 -255
rect 487 -336 887 -289
rect -887 -583 -487 -536
rect -887 -617 -871 -583
rect -503 -617 -487 -583
rect -887 -633 -487 -617
rect -429 -583 -29 -536
rect -429 -617 -413 -583
rect -45 -617 -29 -583
rect -429 -633 -29 -617
rect 29 -583 429 -536
rect 29 -617 45 -583
rect 413 -617 429 -583
rect 29 -633 429 -617
rect 487 -583 887 -536
rect 487 -617 503 -583
rect 871 -617 887 -583
rect 487 -633 887 -617
<< polycont >>
rect -871 583 -503 617
rect -413 583 -45 617
rect 45 583 413 617
rect 503 583 871 617
rect -871 255 -503 289
rect -413 255 -45 289
rect 45 255 413 289
rect 503 255 871 289
rect -871 147 -503 181
rect -413 147 -45 181
rect 45 147 413 181
rect 503 147 871 181
rect -871 -181 -503 -147
rect -413 -181 -45 -147
rect 45 -181 413 -147
rect 503 -181 871 -147
rect -871 -289 -503 -255
rect -413 -289 -45 -255
rect 45 -289 413 -255
rect 503 -289 871 -255
rect -871 -617 -503 -583
rect -413 -617 -45 -583
rect 45 -617 413 -583
rect 503 -617 871 -583
<< locali >>
rect -1047 685 -951 719
rect 951 685 1047 719
rect -1047 623 -1013 685
rect 1013 623 1047 685
rect -887 583 -871 617
rect -503 583 -487 617
rect -429 583 -413 617
rect -45 583 -29 617
rect 29 583 45 617
rect 413 583 429 617
rect 487 583 503 617
rect 871 583 887 617
rect -933 524 -899 540
rect -933 332 -899 348
rect -475 524 -441 540
rect -475 332 -441 348
rect -17 524 17 540
rect -17 332 17 348
rect 441 524 475 540
rect 441 332 475 348
rect 899 524 933 540
rect 899 332 933 348
rect -887 255 -871 289
rect -503 255 -487 289
rect -429 255 -413 289
rect -45 255 -29 289
rect 29 255 45 289
rect 413 255 429 289
rect 487 255 503 289
rect 871 255 887 289
rect -887 147 -871 181
rect -503 147 -487 181
rect -429 147 -413 181
rect -45 147 -29 181
rect 29 147 45 181
rect 413 147 429 181
rect 487 147 503 181
rect 871 147 887 181
rect -933 88 -899 104
rect -933 -104 -899 -88
rect -475 88 -441 104
rect -475 -104 -441 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 441 88 475 104
rect 441 -104 475 -88
rect 899 88 933 104
rect 899 -104 933 -88
rect -887 -181 -871 -147
rect -503 -181 -487 -147
rect -429 -181 -413 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 413 -181 429 -147
rect 487 -181 503 -147
rect 871 -181 887 -147
rect -887 -289 -871 -255
rect -503 -289 -487 -255
rect -429 -289 -413 -255
rect -45 -289 -29 -255
rect 29 -289 45 -255
rect 413 -289 429 -255
rect 487 -289 503 -255
rect 871 -289 887 -255
rect -933 -348 -899 -332
rect -933 -540 -899 -524
rect -475 -348 -441 -332
rect -475 -540 -441 -524
rect -17 -348 17 -332
rect -17 -540 17 -524
rect 441 -348 475 -332
rect 441 -540 475 -524
rect 899 -348 933 -332
rect 899 -540 933 -524
rect -887 -617 -871 -583
rect -503 -617 -487 -583
rect -429 -617 -413 -583
rect -45 -617 -29 -583
rect 29 -617 45 -583
rect 413 -617 429 -583
rect 487 -617 503 -583
rect 871 -617 887 -583
rect -1047 -685 -1013 -623
rect 1013 -685 1047 -623
rect -1047 -719 -951 -685
rect 951 -719 1047 -685
<< viali >>
rect -871 583 -503 617
rect -413 583 -45 617
rect 45 583 413 617
rect 503 583 871 617
rect -933 348 -899 524
rect -475 348 -441 524
rect -17 348 17 524
rect 441 348 475 524
rect 899 348 933 524
rect -871 255 -503 289
rect -413 255 -45 289
rect 45 255 413 289
rect 503 255 871 289
rect -871 147 -503 181
rect -413 147 -45 181
rect 45 147 413 181
rect 503 147 871 181
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect -871 -181 -503 -147
rect -413 -181 -45 -147
rect 45 -181 413 -147
rect 503 -181 871 -147
rect -871 -289 -503 -255
rect -413 -289 -45 -255
rect 45 -289 413 -255
rect 503 -289 871 -255
rect -933 -524 -899 -348
rect -475 -524 -441 -348
rect -17 -524 17 -348
rect 441 -524 475 -348
rect 899 -524 933 -348
rect -871 -617 -503 -583
rect -413 -617 -45 -583
rect 45 -617 413 -583
rect 503 -617 871 -583
<< metal1 >>
rect -883 617 -491 623
rect -883 583 -871 617
rect -503 583 -491 617
rect -883 577 -491 583
rect -425 617 -33 623
rect -425 583 -413 617
rect -45 583 -33 617
rect -425 577 -33 583
rect 33 617 425 623
rect 33 583 45 617
rect 413 583 425 617
rect 33 577 425 583
rect 491 617 883 623
rect 491 583 503 617
rect 871 583 883 617
rect 491 577 883 583
rect -939 524 -893 536
rect -939 348 -933 524
rect -899 348 -893 524
rect -939 336 -893 348
rect -481 524 -435 536
rect -481 348 -475 524
rect -441 348 -435 524
rect -481 336 -435 348
rect -23 524 23 536
rect -23 348 -17 524
rect 17 348 23 524
rect -23 336 23 348
rect 435 524 481 536
rect 435 348 441 524
rect 475 348 481 524
rect 435 336 481 348
rect 893 524 939 536
rect 893 348 899 524
rect 933 348 939 524
rect 893 336 939 348
rect -883 289 -491 295
rect -883 255 -871 289
rect -503 255 -491 289
rect -883 249 -491 255
rect -425 289 -33 295
rect -425 255 -413 289
rect -45 255 -33 289
rect -425 249 -33 255
rect 33 289 425 295
rect 33 255 45 289
rect 413 255 425 289
rect 33 249 425 255
rect 491 289 883 295
rect 491 255 503 289
rect 871 255 883 289
rect 491 249 883 255
rect -883 181 -491 187
rect -883 147 -871 181
rect -503 147 -491 181
rect -883 141 -491 147
rect -425 181 -33 187
rect -425 147 -413 181
rect -45 147 -33 181
rect -425 141 -33 147
rect 33 181 425 187
rect 33 147 45 181
rect 413 147 425 181
rect 33 141 425 147
rect 491 181 883 187
rect 491 147 503 181
rect 871 147 883 181
rect 491 141 883 147
rect -939 88 -893 100
rect -939 -88 -933 88
rect -899 -88 -893 88
rect -939 -100 -893 -88
rect -481 88 -435 100
rect -481 -88 -475 88
rect -441 -88 -435 88
rect -481 -100 -435 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 435 88 481 100
rect 435 -88 441 88
rect 475 -88 481 88
rect 435 -100 481 -88
rect 893 88 939 100
rect 893 -88 899 88
rect 933 -88 939 88
rect 893 -100 939 -88
rect -883 -147 -491 -141
rect -883 -181 -871 -147
rect -503 -181 -491 -147
rect -883 -187 -491 -181
rect -425 -147 -33 -141
rect -425 -181 -413 -147
rect -45 -181 -33 -147
rect -425 -187 -33 -181
rect 33 -147 425 -141
rect 33 -181 45 -147
rect 413 -181 425 -147
rect 33 -187 425 -181
rect 491 -147 883 -141
rect 491 -181 503 -147
rect 871 -181 883 -147
rect 491 -187 883 -181
rect -883 -255 -491 -249
rect -883 -289 -871 -255
rect -503 -289 -491 -255
rect -883 -295 -491 -289
rect -425 -255 -33 -249
rect -425 -289 -413 -255
rect -45 -289 -33 -255
rect -425 -295 -33 -289
rect 33 -255 425 -249
rect 33 -289 45 -255
rect 413 -289 425 -255
rect 33 -295 425 -289
rect 491 -255 883 -249
rect 491 -289 503 -255
rect 871 -289 883 -255
rect 491 -295 883 -289
rect -939 -348 -893 -336
rect -939 -524 -933 -348
rect -899 -524 -893 -348
rect -939 -536 -893 -524
rect -481 -348 -435 -336
rect -481 -524 -475 -348
rect -441 -524 -435 -348
rect -481 -536 -435 -524
rect -23 -348 23 -336
rect -23 -524 -17 -348
rect 17 -524 23 -348
rect -23 -536 23 -524
rect 435 -348 481 -336
rect 435 -524 441 -348
rect 475 -524 481 -348
rect 435 -536 481 -524
rect 893 -348 939 -336
rect 893 -524 899 -348
rect 933 -524 939 -348
rect 893 -536 939 -524
rect -883 -583 -491 -577
rect -883 -617 -871 -583
rect -503 -617 -491 -583
rect -883 -623 -491 -617
rect -425 -583 -33 -577
rect -425 -617 -413 -583
rect -45 -617 -33 -583
rect -425 -623 -33 -617
rect 33 -583 425 -577
rect 33 -617 45 -583
rect 413 -617 425 -583
rect 33 -623 425 -617
rect 491 -583 883 -577
rect 491 -617 503 -583
rect 871 -617 883 -583
rect 491 -623 883 -617
<< properties >>
string FIXED_BBOX -1030 -702 1030 702
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 2 m 3 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
