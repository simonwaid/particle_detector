magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< error_p >>
rect -173 272 -115 278
rect 19 272 77 278
rect 211 272 269 278
rect -173 238 -161 272
rect 19 238 31 272
rect 211 238 223 272
rect -173 232 -115 238
rect 19 232 77 238
rect 211 232 269 238
rect -269 -238 -211 -232
rect -77 -238 -19 -232
rect 115 -238 173 -232
rect -269 -272 -257 -238
rect -77 -272 -65 -238
rect 115 -272 127 -238
rect -269 -278 -211 -272
rect -77 -278 -19 -272
rect 115 -278 173 -272
<< pwell >>
rect -455 -410 455 410
<< nmoslvt >>
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
<< ndiff >>
rect -317 188 -255 200
rect -317 -188 -305 188
rect -271 -188 -255 188
rect -317 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 317 200
rect 255 -188 271 188
rect 305 -188 317 188
rect 255 -200 317 -188
<< ndiffc >>
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
<< psubdiff >>
rect -419 340 -323 374
rect 323 340 419 374
rect -419 278 -385 340
rect 385 278 419 340
rect -419 -340 -385 -278
rect 385 -340 419 -278
rect -419 -374 -323 -340
rect 323 -374 419 -340
<< psubdiffcont >>
rect -323 340 323 374
rect -419 -278 -385 278
rect 385 -278 419 278
rect -323 -374 323 -340
<< poly >>
rect -177 272 -111 288
rect -177 238 -161 272
rect -127 238 -111 272
rect -255 200 -225 226
rect -177 222 -111 238
rect 15 272 81 288
rect 15 238 31 272
rect 65 238 81 272
rect -159 200 -129 222
rect -63 200 -33 226
rect 15 222 81 238
rect 207 272 273 288
rect 207 238 223 272
rect 257 238 273 272
rect 33 200 63 222
rect 129 200 159 226
rect 207 222 273 238
rect 225 200 255 222
rect -255 -222 -225 -200
rect -273 -238 -207 -222
rect -159 -226 -129 -200
rect -63 -222 -33 -200
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -273 -288 -207 -272
rect -81 -238 -15 -222
rect 33 -226 63 -200
rect 129 -222 159 -200
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect -81 -288 -15 -272
rect 111 -238 177 -222
rect 225 -226 255 -200
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 111 -288 177 -272
<< polycont >>
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
<< locali >>
rect -419 340 -323 374
rect 323 340 419 374
rect -419 278 -385 340
rect 385 278 419 340
rect -177 238 -161 272
rect -127 238 -111 272
rect 15 238 31 272
rect 65 238 81 272
rect 207 238 223 272
rect 257 238 273 272
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect 111 -272 127 -238
rect 161 -272 177 -238
rect -419 -340 -385 -278
rect 385 -340 419 -278
rect -419 -374 -323 -340
rect 323 -374 419 -340
<< viali >>
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
<< metal1 >>
rect -173 272 -115 278
rect -173 238 -161 272
rect -127 238 -115 272
rect -173 232 -115 238
rect 19 272 77 278
rect 19 238 31 272
rect 65 238 77 272
rect 19 232 77 238
rect 211 272 269 278
rect 211 238 223 272
rect 257 238 269 272
rect 211 232 269 238
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect -269 -238 -211 -232
rect -269 -272 -257 -238
rect -223 -272 -211 -238
rect -269 -278 -211 -272
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -31 -272 -19 -238
rect -77 -278 -19 -272
rect 115 -238 173 -232
rect 115 -272 127 -238
rect 161 -272 173 -238
rect 115 -278 173 -272
<< properties >>
string FIXED_BBOX -402 -357 402 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
