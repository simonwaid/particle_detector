magic
tech sky130A
magscale 1 2
timestamp 1645541123
<< error_p >>
rect -6670 591 -6210 618
rect -5750 591 -5290 618
rect -4830 591 -4370 618
rect -3910 591 -3450 618
rect -2990 591 -2530 618
rect -2070 591 -1610 618
rect -6670 -618 -6210 -591
rect -5750 -618 -5290 -591
rect -4830 -618 -4370 -591
rect -3910 -618 -3450 -591
rect -2990 -618 -2530 -591
rect -2070 -618 -1610 -591
<< nwell >>
rect -6773 -591 -6107 591
rect -5853 -591 -5187 591
rect -4933 -591 -4267 591
rect -4013 -591 -3347 591
rect -3093 -591 -2427 591
rect -2173 -591 -1507 591
rect -1253 -591 -587 591
rect -333 -591 333 591
rect 587 -591 1253 591
rect 1507 -591 2173 591
rect 2427 -591 3093 591
rect 3347 -591 4013 591
rect 4267 -591 4933 591
rect 5187 -591 5853 591
rect 6107 -591 6773 591
<< pwell >>
rect -6883 591 6883 701
rect -6883 -591 -6773 591
rect -6107 -591 -5853 591
rect -5187 -591 -4933 591
rect -4267 -591 -4013 591
rect -3347 -591 -3093 591
rect -2427 -591 -2173 591
rect -1507 -591 -1253 591
rect -587 -591 -333 591
rect 333 -591 587 591
rect 1253 -591 1507 591
rect 2173 -591 2427 591
rect 3093 -591 3347 591
rect 4013 -591 4267 591
rect 4933 -591 5187 591
rect 5853 -591 6107 591
rect 6773 -591 6883 591
rect -6883 -701 6883 -591
<< varactor >>
rect -6640 -500 -6240 500
rect -5720 -500 -5320 500
rect -4800 -500 -4400 500
rect -3880 -500 -3480 500
rect -2960 -500 -2560 500
rect -2040 -500 -1640 500
rect -1120 -500 -720 500
rect -200 -500 200 500
rect 720 -500 1120 500
rect 1640 -500 2040 500
rect 2560 -500 2960 500
rect 3480 -500 3880 500
rect 4400 -500 4800 500
rect 5320 -500 5720 500
rect 6240 -500 6640 500
<< psubdiff >>
rect -6847 631 -6751 665
rect 6751 631 6847 665
rect -6847 569 -6813 631
rect 6813 569 6847 631
rect -6847 -631 -6813 -569
rect 6813 -631 6847 -569
rect -6847 -665 -6751 -631
rect 6751 -665 6847 -631
<< nsubdiff >>
rect -6737 476 -6640 500
rect -6737 -476 -6725 476
rect -6691 -476 -6640 476
rect -6737 -500 -6640 -476
rect -6240 476 -6143 500
rect -6240 -476 -6189 476
rect -6155 -476 -6143 476
rect -6240 -500 -6143 -476
rect -5817 476 -5720 500
rect -5817 -476 -5805 476
rect -5771 -476 -5720 476
rect -5817 -500 -5720 -476
rect -5320 476 -5223 500
rect -5320 -476 -5269 476
rect -5235 -476 -5223 476
rect -5320 -500 -5223 -476
rect -4897 476 -4800 500
rect -4897 -476 -4885 476
rect -4851 -476 -4800 476
rect -4897 -500 -4800 -476
rect -4400 476 -4303 500
rect -4400 -476 -4349 476
rect -4315 -476 -4303 476
rect -4400 -500 -4303 -476
rect -3977 476 -3880 500
rect -3977 -476 -3965 476
rect -3931 -476 -3880 476
rect -3977 -500 -3880 -476
rect -3480 476 -3383 500
rect -3480 -476 -3429 476
rect -3395 -476 -3383 476
rect -3480 -500 -3383 -476
rect -3057 476 -2960 500
rect -3057 -476 -3045 476
rect -3011 -476 -2960 476
rect -3057 -500 -2960 -476
rect -2560 476 -2463 500
rect -2560 -476 -2509 476
rect -2475 -476 -2463 476
rect -2560 -500 -2463 -476
rect -2137 476 -2040 500
rect -2137 -476 -2125 476
rect -2091 -476 -2040 476
rect -2137 -500 -2040 -476
rect -1640 476 -1543 500
rect -1640 -476 -1589 476
rect -1555 -476 -1543 476
rect -1640 -500 -1543 -476
rect -1217 476 -1120 500
rect -1217 -476 -1205 476
rect -1171 -476 -1120 476
rect -1217 -500 -1120 -476
rect -720 476 -623 500
rect -720 -476 -669 476
rect -635 -476 -623 476
rect -720 -500 -623 -476
rect -297 476 -200 500
rect -297 -476 -285 476
rect -251 -476 -200 476
rect -297 -500 -200 -476
rect 200 476 297 500
rect 200 -476 251 476
rect 285 -476 297 476
rect 200 -500 297 -476
rect 623 476 720 500
rect 623 -476 635 476
rect 669 -476 720 476
rect 623 -500 720 -476
rect 1120 476 1217 500
rect 1120 -476 1171 476
rect 1205 -476 1217 476
rect 1120 -500 1217 -476
rect 1543 476 1640 500
rect 1543 -476 1555 476
rect 1589 -476 1640 476
rect 1543 -500 1640 -476
rect 2040 476 2137 500
rect 2040 -476 2091 476
rect 2125 -476 2137 476
rect 2040 -500 2137 -476
rect 2463 476 2560 500
rect 2463 -476 2475 476
rect 2509 -476 2560 476
rect 2463 -500 2560 -476
rect 2960 476 3057 500
rect 2960 -476 3011 476
rect 3045 -476 3057 476
rect 2960 -500 3057 -476
rect 3383 476 3480 500
rect 3383 -476 3395 476
rect 3429 -476 3480 476
rect 3383 -500 3480 -476
rect 3880 476 3977 500
rect 3880 -476 3931 476
rect 3965 -476 3977 476
rect 3880 -500 3977 -476
rect 4303 476 4400 500
rect 4303 -476 4315 476
rect 4349 -476 4400 476
rect 4303 -500 4400 -476
rect 4800 476 4897 500
rect 4800 -476 4851 476
rect 4885 -476 4897 476
rect 4800 -500 4897 -476
rect 5223 476 5320 500
rect 5223 -476 5235 476
rect 5269 -476 5320 476
rect 5223 -500 5320 -476
rect 5720 476 5817 500
rect 5720 -476 5771 476
rect 5805 -476 5817 476
rect 5720 -500 5817 -476
rect 6143 476 6240 500
rect 6143 -476 6155 476
rect 6189 -476 6240 476
rect 6143 -500 6240 -476
rect 6640 476 6737 500
rect 6640 -476 6691 476
rect 6725 -476 6737 476
rect 6640 -500 6737 -476
<< psubdiffcont >>
rect -6751 631 6751 665
rect -6847 -569 -6813 569
rect 6813 -569 6847 569
rect -6751 -665 6751 -631
<< nsubdiffcont >>
rect -6725 -476 -6691 476
rect -6189 -476 -6155 476
rect -5805 -476 -5771 476
rect -5269 -476 -5235 476
rect -4885 -476 -4851 476
rect -4349 -476 -4315 476
rect -3965 -476 -3931 476
rect -3429 -476 -3395 476
rect -3045 -476 -3011 476
rect -2509 -476 -2475 476
rect -2125 -476 -2091 476
rect -1589 -476 -1555 476
rect -1205 -476 -1171 476
rect -669 -476 -635 476
rect -285 -476 -251 476
rect 251 -476 285 476
rect 635 -476 669 476
rect 1171 -476 1205 476
rect 1555 -476 1589 476
rect 2091 -476 2125 476
rect 2475 -476 2509 476
rect 3011 -476 3045 476
rect 3395 -476 3429 476
rect 3931 -476 3965 476
rect 4315 -476 4349 476
rect 4851 -476 4885 476
rect 5235 -476 5269 476
rect 5771 -476 5805 476
rect 6155 -476 6189 476
rect 6691 -476 6725 476
<< poly >>
rect -6640 572 -6240 588
rect -6640 538 -6624 572
rect -6256 538 -6240 572
rect -6640 500 -6240 538
rect -5720 572 -5320 588
rect -5720 538 -5704 572
rect -5336 538 -5320 572
rect -5720 500 -5320 538
rect -4800 572 -4400 588
rect -4800 538 -4784 572
rect -4416 538 -4400 572
rect -4800 500 -4400 538
rect -3880 572 -3480 588
rect -3880 538 -3864 572
rect -3496 538 -3480 572
rect -3880 500 -3480 538
rect -2960 572 -2560 588
rect -2960 538 -2944 572
rect -2576 538 -2560 572
rect -2960 500 -2560 538
rect -2040 572 -1640 588
rect -2040 538 -2024 572
rect -1656 538 -1640 572
rect -2040 500 -1640 538
rect -1120 572 -720 588
rect -1120 538 -1104 572
rect -736 538 -720 572
rect -1120 500 -720 538
rect -200 572 200 588
rect -200 538 -184 572
rect 184 538 200 572
rect -200 500 200 538
rect 720 572 1120 588
rect 720 538 736 572
rect 1104 538 1120 572
rect 720 500 1120 538
rect 1640 572 2040 588
rect 1640 538 1656 572
rect 2024 538 2040 572
rect 1640 500 2040 538
rect 2560 572 2960 588
rect 2560 538 2576 572
rect 2944 538 2960 572
rect 2560 500 2960 538
rect 3480 572 3880 588
rect 3480 538 3496 572
rect 3864 538 3880 572
rect 3480 500 3880 538
rect 4400 572 4800 588
rect 4400 538 4416 572
rect 4784 538 4800 572
rect 4400 500 4800 538
rect 5320 572 5720 588
rect 5320 538 5336 572
rect 5704 538 5720 572
rect 5320 500 5720 538
rect 6240 572 6640 588
rect 6240 538 6256 572
rect 6624 538 6640 572
rect 6240 500 6640 538
rect -6640 -538 -6240 -500
rect -6640 -572 -6624 -538
rect -6256 -572 -6240 -538
rect -6640 -588 -6240 -572
rect -5720 -538 -5320 -500
rect -5720 -572 -5704 -538
rect -5336 -572 -5320 -538
rect -5720 -588 -5320 -572
rect -4800 -538 -4400 -500
rect -4800 -572 -4784 -538
rect -4416 -572 -4400 -538
rect -4800 -588 -4400 -572
rect -3880 -538 -3480 -500
rect -3880 -572 -3864 -538
rect -3496 -572 -3480 -538
rect -3880 -588 -3480 -572
rect -2960 -538 -2560 -500
rect -2960 -572 -2944 -538
rect -2576 -572 -2560 -538
rect -2960 -588 -2560 -572
rect -2040 -538 -1640 -500
rect -2040 -572 -2024 -538
rect -1656 -572 -1640 -538
rect -2040 -588 -1640 -572
rect -1120 -538 -720 -500
rect -1120 -572 -1104 -538
rect -736 -572 -720 -538
rect -1120 -588 -720 -572
rect -200 -538 200 -500
rect -200 -572 -184 -538
rect 184 -572 200 -538
rect -200 -588 200 -572
rect 720 -538 1120 -500
rect 720 -572 736 -538
rect 1104 -572 1120 -538
rect 720 -588 1120 -572
rect 1640 -538 2040 -500
rect 1640 -572 1656 -538
rect 2024 -572 2040 -538
rect 1640 -588 2040 -572
rect 2560 -538 2960 -500
rect 2560 -572 2576 -538
rect 2944 -572 2960 -538
rect 2560 -588 2960 -572
rect 3480 -538 3880 -500
rect 3480 -572 3496 -538
rect 3864 -572 3880 -538
rect 3480 -588 3880 -572
rect 4400 -538 4800 -500
rect 4400 -572 4416 -538
rect 4784 -572 4800 -538
rect 4400 -588 4800 -572
rect 5320 -538 5720 -500
rect 5320 -572 5336 -538
rect 5704 -572 5720 -538
rect 5320 -588 5720 -572
rect 6240 -538 6640 -500
rect 6240 -572 6256 -538
rect 6624 -572 6640 -538
rect 6240 -588 6640 -572
<< polycont >>
rect -6624 538 -6256 572
rect -5704 538 -5336 572
rect -4784 538 -4416 572
rect -3864 538 -3496 572
rect -2944 538 -2576 572
rect -2024 538 -1656 572
rect -1104 538 -736 572
rect -184 538 184 572
rect 736 538 1104 572
rect 1656 538 2024 572
rect 2576 538 2944 572
rect 3496 538 3864 572
rect 4416 538 4784 572
rect 5336 538 5704 572
rect 6256 538 6624 572
rect -6624 -572 -6256 -538
rect -5704 -572 -5336 -538
rect -4784 -572 -4416 -538
rect -3864 -572 -3496 -538
rect -2944 -572 -2576 -538
rect -2024 -572 -1656 -538
rect -1104 -572 -736 -538
rect -184 -572 184 -538
rect 736 -572 1104 -538
rect 1656 -572 2024 -538
rect 2576 -572 2944 -538
rect 3496 -572 3864 -538
rect 4416 -572 4784 -538
rect 5336 -572 5704 -538
rect 6256 -572 6624 -538
<< locali >>
rect -6847 631 -6751 665
rect 6751 631 6847 665
rect -6847 569 -6813 631
rect -6640 538 -6624 572
rect -6256 538 -6240 572
rect -5720 538 -5704 572
rect -5336 538 -5320 572
rect -4800 538 -4784 572
rect -4416 538 -4400 572
rect -3880 538 -3864 572
rect -3496 538 -3480 572
rect -2960 538 -2944 572
rect -2576 538 -2560 572
rect -2040 538 -2024 572
rect -1656 538 -1640 572
rect -1120 538 -1104 572
rect -736 538 -720 572
rect -200 538 -184 572
rect 184 538 200 572
rect 720 538 736 572
rect 1104 538 1120 572
rect 1640 538 1656 572
rect 2024 538 2040 572
rect 2560 538 2576 572
rect 2944 538 2960 572
rect 3480 538 3496 572
rect 3864 538 3880 572
rect 4400 538 4416 572
rect 4784 538 4800 572
rect 5320 538 5336 572
rect 5704 538 5720 572
rect 6240 538 6256 572
rect 6624 538 6640 572
rect 6813 569 6847 631
rect -6725 476 -6691 492
rect -6725 -492 -6691 -476
rect -6189 476 -6155 492
rect -6189 -492 -6155 -476
rect -5805 476 -5771 492
rect -5805 -492 -5771 -476
rect -5269 476 -5235 492
rect -5269 -492 -5235 -476
rect -4885 476 -4851 492
rect -4885 -492 -4851 -476
rect -4349 476 -4315 492
rect -4349 -492 -4315 -476
rect -3965 476 -3931 492
rect -3965 -492 -3931 -476
rect -3429 476 -3395 492
rect -3429 -492 -3395 -476
rect -3045 476 -3011 492
rect -3045 -492 -3011 -476
rect -2509 476 -2475 492
rect -2509 -492 -2475 -476
rect -2125 476 -2091 492
rect -2125 -492 -2091 -476
rect -1589 476 -1555 492
rect -1589 -492 -1555 -476
rect -1205 476 -1171 492
rect -1205 -492 -1171 -476
rect -669 476 -635 492
rect -669 -492 -635 -476
rect -285 476 -251 492
rect -285 -492 -251 -476
rect 251 476 285 492
rect 251 -492 285 -476
rect 635 476 669 492
rect 635 -492 669 -476
rect 1171 476 1205 492
rect 1171 -492 1205 -476
rect 1555 476 1589 492
rect 1555 -492 1589 -476
rect 2091 476 2125 492
rect 2091 -492 2125 -476
rect 2475 476 2509 492
rect 2475 -492 2509 -476
rect 3011 476 3045 492
rect 3011 -492 3045 -476
rect 3395 476 3429 492
rect 3395 -492 3429 -476
rect 3931 476 3965 492
rect 3931 -492 3965 -476
rect 4315 476 4349 492
rect 4315 -492 4349 -476
rect 4851 476 4885 492
rect 4851 -492 4885 -476
rect 5235 476 5269 492
rect 5235 -492 5269 -476
rect 5771 476 5805 492
rect 5771 -492 5805 -476
rect 6155 476 6189 492
rect 6155 -492 6189 -476
rect 6691 476 6725 492
rect 6691 -492 6725 -476
rect -6847 -631 -6813 -569
rect -6640 -572 -6624 -538
rect -6256 -572 -6240 -538
rect -5720 -572 -5704 -538
rect -5336 -572 -5320 -538
rect -4800 -572 -4784 -538
rect -4416 -572 -4400 -538
rect -3880 -572 -3864 -538
rect -3496 -572 -3480 -538
rect -2960 -572 -2944 -538
rect -2576 -572 -2560 -538
rect -2040 -572 -2024 -538
rect -1656 -572 -1640 -538
rect -1120 -572 -1104 -538
rect -736 -572 -720 -538
rect -200 -572 -184 -538
rect 184 -572 200 -538
rect 720 -572 736 -538
rect 1104 -572 1120 -538
rect 1640 -572 1656 -538
rect 2024 -572 2040 -538
rect 2560 -572 2576 -538
rect 2944 -572 2960 -538
rect 3480 -572 3496 -538
rect 3864 -572 3880 -538
rect 4400 -572 4416 -538
rect 4784 -572 4800 -538
rect 5320 -572 5336 -538
rect 5704 -572 5720 -538
rect 6240 -572 6256 -538
rect 6624 -572 6640 -538
rect 6813 -631 6847 -569
rect -6847 -665 -6751 -631
rect 6751 -665 6847 -631
<< viali >>
rect -6624 538 -6256 572
rect -5704 538 -5336 572
rect -4784 538 -4416 572
rect -3864 538 -3496 572
rect -2944 538 -2576 572
rect -2024 538 -1656 572
rect -1104 538 -736 572
rect -184 538 184 572
rect 736 538 1104 572
rect 1656 538 2024 572
rect 2576 538 2944 572
rect 3496 538 3864 572
rect 4416 538 4784 572
rect 5336 538 5704 572
rect 6256 538 6624 572
rect -6725 -476 -6691 476
rect -6189 -476 -6155 476
rect -5805 -476 -5771 476
rect -5269 -476 -5235 476
rect -4885 -476 -4851 476
rect -4349 -476 -4315 476
rect -3965 -476 -3931 476
rect -3429 -476 -3395 476
rect -3045 -476 -3011 476
rect -2509 -476 -2475 476
rect -2125 -476 -2091 476
rect -1589 -476 -1555 476
rect -1205 -476 -1171 476
rect -669 -476 -635 476
rect -285 -476 -251 476
rect 251 -476 285 476
rect 635 -476 669 476
rect 1171 -476 1205 476
rect 1555 -476 1589 476
rect 2091 -476 2125 476
rect 2475 -476 2509 476
rect 3011 -476 3045 476
rect 3395 -476 3429 476
rect 3931 -476 3965 476
rect 4315 -476 4349 476
rect 4851 -476 4885 476
rect 5235 -476 5269 476
rect 5771 -476 5805 476
rect 6155 -476 6189 476
rect 6691 -476 6725 476
rect -6624 -572 -6256 -538
rect -5704 -572 -5336 -538
rect -4784 -572 -4416 -538
rect -3864 -572 -3496 -538
rect -2944 -572 -2576 -538
rect -2024 -572 -1656 -538
rect -1104 -572 -736 -538
rect -184 -572 184 -538
rect 736 -572 1104 -538
rect 1656 -572 2024 -538
rect 2576 -572 2944 -538
rect 3496 -572 3864 -538
rect 4416 -572 4784 -538
rect 5336 -572 5704 -538
rect 6256 -572 6624 -538
<< metal1 >>
rect -6636 572 -6244 578
rect -6636 538 -6624 572
rect -6256 538 -6244 572
rect -6636 532 -6244 538
rect -5716 572 -5324 578
rect -5716 538 -5704 572
rect -5336 538 -5324 572
rect -5716 532 -5324 538
rect -4796 572 -4404 578
rect -4796 538 -4784 572
rect -4416 538 -4404 572
rect -4796 532 -4404 538
rect -3876 572 -3484 578
rect -3876 538 -3864 572
rect -3496 538 -3484 572
rect -3876 532 -3484 538
rect -2956 572 -2564 578
rect -2956 538 -2944 572
rect -2576 538 -2564 572
rect -2956 532 -2564 538
rect -2036 572 -1644 578
rect -2036 538 -2024 572
rect -1656 538 -1644 572
rect -2036 532 -1644 538
rect -1116 572 -724 578
rect -1116 538 -1104 572
rect -736 538 -724 572
rect -1116 532 -724 538
rect -196 572 196 578
rect -196 538 -184 572
rect 184 538 196 572
rect -196 532 196 538
rect 724 572 1116 578
rect 724 538 736 572
rect 1104 538 1116 572
rect 724 532 1116 538
rect 1644 572 2036 578
rect 1644 538 1656 572
rect 2024 538 2036 572
rect 1644 532 2036 538
rect 2564 572 2956 578
rect 2564 538 2576 572
rect 2944 538 2956 572
rect 2564 532 2956 538
rect 3484 572 3876 578
rect 3484 538 3496 572
rect 3864 538 3876 572
rect 3484 532 3876 538
rect 4404 572 4796 578
rect 4404 538 4416 572
rect 4784 538 4796 572
rect 4404 532 4796 538
rect 5324 572 5716 578
rect 5324 538 5336 572
rect 5704 538 5716 572
rect 5324 532 5716 538
rect 6244 572 6636 578
rect 6244 538 6256 572
rect 6624 538 6636 572
rect 6244 532 6636 538
rect -6731 476 -6685 488
rect -6731 -476 -6725 476
rect -6691 -476 -6685 476
rect -6731 -488 -6685 -476
rect -6195 476 -6149 488
rect -6195 -476 -6189 476
rect -6155 -476 -6149 476
rect -6195 -488 -6149 -476
rect -5811 476 -5765 488
rect -5811 -476 -5805 476
rect -5771 -476 -5765 476
rect -5811 -488 -5765 -476
rect -5275 476 -5229 488
rect -5275 -476 -5269 476
rect -5235 -476 -5229 476
rect -5275 -488 -5229 -476
rect -4891 476 -4845 488
rect -4891 -476 -4885 476
rect -4851 -476 -4845 476
rect -4891 -488 -4845 -476
rect -4355 476 -4309 488
rect -4355 -476 -4349 476
rect -4315 -476 -4309 476
rect -4355 -488 -4309 -476
rect -3971 476 -3925 488
rect -3971 -476 -3965 476
rect -3931 -476 -3925 476
rect -3971 -488 -3925 -476
rect -3435 476 -3389 488
rect -3435 -476 -3429 476
rect -3395 -476 -3389 476
rect -3435 -488 -3389 -476
rect -3051 476 -3005 488
rect -3051 -476 -3045 476
rect -3011 -476 -3005 476
rect -3051 -488 -3005 -476
rect -2515 476 -2469 488
rect -2515 -476 -2509 476
rect -2475 -476 -2469 476
rect -2515 -488 -2469 -476
rect -2131 476 -2085 488
rect -2131 -476 -2125 476
rect -2091 -476 -2085 476
rect -2131 -488 -2085 -476
rect -1595 476 -1549 488
rect -1595 -476 -1589 476
rect -1555 -476 -1549 476
rect -1595 -488 -1549 -476
rect -1211 476 -1165 488
rect -1211 -476 -1205 476
rect -1171 -476 -1165 476
rect -1211 -488 -1165 -476
rect -675 476 -629 488
rect -675 -476 -669 476
rect -635 -476 -629 476
rect -675 -488 -629 -476
rect -291 476 -245 488
rect -291 -476 -285 476
rect -251 -476 -245 476
rect -291 -488 -245 -476
rect 245 476 291 488
rect 245 -476 251 476
rect 285 -476 291 476
rect 245 -488 291 -476
rect 629 476 675 488
rect 629 -476 635 476
rect 669 -476 675 476
rect 629 -488 675 -476
rect 1165 476 1211 488
rect 1165 -476 1171 476
rect 1205 -476 1211 476
rect 1165 -488 1211 -476
rect 1549 476 1595 488
rect 1549 -476 1555 476
rect 1589 -476 1595 476
rect 1549 -488 1595 -476
rect 2085 476 2131 488
rect 2085 -476 2091 476
rect 2125 -476 2131 476
rect 2085 -488 2131 -476
rect 2469 476 2515 488
rect 2469 -476 2475 476
rect 2509 -476 2515 476
rect 2469 -488 2515 -476
rect 3005 476 3051 488
rect 3005 -476 3011 476
rect 3045 -476 3051 476
rect 3005 -488 3051 -476
rect 3389 476 3435 488
rect 3389 -476 3395 476
rect 3429 -476 3435 476
rect 3389 -488 3435 -476
rect 3925 476 3971 488
rect 3925 -476 3931 476
rect 3965 -476 3971 476
rect 3925 -488 3971 -476
rect 4309 476 4355 488
rect 4309 -476 4315 476
rect 4349 -476 4355 476
rect 4309 -488 4355 -476
rect 4845 476 4891 488
rect 4845 -476 4851 476
rect 4885 -476 4891 476
rect 4845 -488 4891 -476
rect 5229 476 5275 488
rect 5229 -476 5235 476
rect 5269 -476 5275 476
rect 5229 -488 5275 -476
rect 5765 476 5811 488
rect 5765 -476 5771 476
rect 5805 -476 5811 476
rect 5765 -488 5811 -476
rect 6149 476 6195 488
rect 6149 -476 6155 476
rect 6189 -476 6195 476
rect 6149 -488 6195 -476
rect 6685 476 6731 488
rect 6685 -476 6691 476
rect 6725 -476 6731 476
rect 6685 -488 6731 -476
rect -6636 -538 -6244 -532
rect -6636 -572 -6624 -538
rect -6256 -572 -6244 -538
rect -6636 -578 -6244 -572
rect -5716 -538 -5324 -532
rect -5716 -572 -5704 -538
rect -5336 -572 -5324 -538
rect -5716 -578 -5324 -572
rect -4796 -538 -4404 -532
rect -4796 -572 -4784 -538
rect -4416 -572 -4404 -538
rect -4796 -578 -4404 -572
rect -3876 -538 -3484 -532
rect -3876 -572 -3864 -538
rect -3496 -572 -3484 -538
rect -3876 -578 -3484 -572
rect -2956 -538 -2564 -532
rect -2956 -572 -2944 -538
rect -2576 -572 -2564 -538
rect -2956 -578 -2564 -572
rect -2036 -538 -1644 -532
rect -2036 -572 -2024 -538
rect -1656 -572 -1644 -538
rect -2036 -578 -1644 -572
rect -1116 -538 -724 -532
rect -1116 -572 -1104 -538
rect -736 -572 -724 -538
rect -1116 -578 -724 -572
rect -196 -538 196 -532
rect -196 -572 -184 -538
rect 184 -572 196 -538
rect -196 -578 196 -572
rect 724 -538 1116 -532
rect 724 -572 736 -538
rect 1104 -572 1116 -538
rect 724 -578 1116 -572
rect 1644 -538 2036 -532
rect 1644 -572 1656 -538
rect 2024 -572 2036 -538
rect 1644 -578 2036 -572
rect 2564 -538 2956 -532
rect 2564 -572 2576 -538
rect 2944 -572 2956 -538
rect 2564 -578 2956 -572
rect 3484 -538 3876 -532
rect 3484 -572 3496 -538
rect 3864 -572 3876 -538
rect 3484 -578 3876 -572
rect 4404 -538 4796 -532
rect 4404 -572 4416 -538
rect 4784 -572 4796 -538
rect 4404 -578 4796 -572
rect 5324 -538 5716 -532
rect 5324 -572 5336 -538
rect 5704 -572 5716 -538
rect 5324 -578 5716 -572
rect 6244 -538 6636 -532
rect 6244 -572 6256 -538
rect 6624 -572 6636 -538
rect 6244 -578 6636 -572
<< properties >>
string FIXED_BBOX -6830 -648 6830 648
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 5 l 2 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
