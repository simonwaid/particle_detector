magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< nwell >>
rect 1482 3720 1644 3786
rect 1992 3720 2154 3786
rect 3192 3720 3546 3786
rect 3892 3720 4246 3786
rect 4592 3720 4754 3786
rect 5102 3720 5456 3786
rect 5802 3720 6156 3786
rect 1500 3706 1530 3720
rect 2010 3708 2040 3720
rect 3210 3706 3240 3720
rect 3402 3702 3432 3720
rect 3910 3704 3940 3720
rect 4102 3698 4132 3720
rect 4610 3704 4640 3720
rect 5120 3708 5150 3720
rect 5312 3706 5342 3720
rect 5820 3700 5850 3720
rect 6012 3702 6042 3720
rect 1596 3258 1626 3270
rect 2106 3258 2136 3276
rect 3306 3258 3336 3280
rect 3498 3258 3528 3278
rect 4006 3258 4036 3280
rect 4198 3258 4228 3278
rect 4706 3258 4736 3272
rect 5216 3258 5246 3274
rect 5408 3258 5438 3276
rect 5916 3258 5946 3284
rect 6108 3258 6138 3284
rect 1546 3248 1644 3258
rect 1482 3202 1644 3248
rect 1546 3192 1644 3202
rect 1992 3192 2154 3258
rect 3192 3192 3546 3258
rect 3892 3192 4246 3258
rect 4592 3192 4754 3258
rect 5102 3192 5456 3258
rect 5802 3192 6156 3258
<< pwell >>
rect 1482 2938 1584 2948
rect 1482 2892 1644 2938
rect 1482 2882 1584 2892
rect 1992 2882 2154 2948
rect 3302 2882 3560 2948
rect 3912 2882 4170 2948
rect 5102 2882 5264 2948
rect 5802 2882 5964 2948
rect 1540 2428 1644 2438
rect 2054 2428 2154 2438
rect 1482 2382 1644 2428
rect 1992 2382 2154 2428
rect 1540 2372 1644 2382
rect 2054 2372 2154 2382
rect 3302 2372 3560 2438
rect 3912 2372 4170 2438
rect 5102 2372 5264 2438
rect 5802 2372 5964 2438
<< poly >>
rect 1482 3770 1644 3786
rect 1482 3736 1498 3770
rect 1532 3736 1644 3770
rect 1482 3720 1644 3736
rect 1992 3770 2154 3786
rect 1992 3736 2008 3770
rect 2042 3736 2154 3770
rect 1992 3720 2154 3736
rect 3192 3770 3546 3786
rect 3192 3736 3208 3770
rect 3242 3736 3400 3770
rect 3434 3736 3546 3770
rect 3192 3720 3546 3736
rect 3892 3770 4246 3786
rect 3892 3736 3908 3770
rect 3942 3736 4100 3770
rect 4134 3736 4246 3770
rect 3892 3720 4246 3736
rect 4592 3770 4754 3786
rect 4592 3736 4608 3770
rect 4642 3736 4754 3770
rect 4592 3720 4754 3736
rect 5102 3770 5456 3786
rect 5102 3736 5118 3770
rect 5152 3736 5310 3770
rect 5344 3736 5456 3770
rect 5102 3720 5456 3736
rect 5802 3770 6156 3786
rect 5802 3736 5818 3770
rect 5852 3736 6010 3770
rect 6044 3736 6156 3770
rect 5802 3720 6156 3736
rect 1500 3706 1530 3720
rect 2010 3708 2040 3720
rect 3210 3706 3240 3720
rect 3402 3702 3432 3720
rect 3910 3704 3940 3720
rect 4102 3698 4132 3720
rect 4610 3704 4640 3720
rect 5120 3708 5150 3720
rect 5312 3706 5342 3720
rect 5820 3700 5850 3720
rect 6012 3702 6042 3720
rect 1596 3258 1626 3270
rect 2106 3258 2136 3276
rect 3306 3258 3336 3280
rect 3498 3258 3528 3278
rect 4006 3258 4036 3280
rect 4198 3258 4228 3278
rect 4706 3258 4736 3272
rect 5216 3258 5246 3274
rect 5408 3258 5438 3276
rect 5916 3258 5946 3284
rect 6108 3258 6138 3284
rect 1546 3248 1644 3258
rect 1482 3242 1644 3248
rect 1482 3208 1594 3242
rect 1628 3208 1644 3242
rect 1482 3202 1644 3208
rect 1546 3192 1644 3202
rect 1992 3242 2154 3258
rect 1992 3208 2104 3242
rect 2138 3208 2154 3242
rect 1992 3192 2154 3208
rect 3192 3242 3546 3258
rect 3192 3208 3304 3242
rect 3338 3208 3496 3242
rect 3530 3208 3546 3242
rect 3192 3192 3546 3208
rect 3892 3242 4246 3258
rect 3892 3208 4004 3242
rect 4038 3208 4196 3242
rect 4230 3208 4246 3242
rect 3892 3192 4246 3208
rect 4592 3242 4754 3258
rect 4592 3208 4704 3242
rect 4738 3208 4754 3242
rect 4592 3192 4754 3208
rect 5102 3242 5456 3258
rect 5102 3208 5214 3242
rect 5248 3208 5406 3242
rect 5440 3208 5456 3242
rect 5102 3192 5456 3208
rect 5802 3242 6156 3258
rect 5802 3208 5914 3242
rect 5948 3208 6106 3242
rect 6140 3208 6156 3242
rect 5802 3192 6156 3208
rect 1482 2938 1584 2948
rect 1482 2932 1644 2938
rect 1482 2898 1498 2932
rect 1532 2898 1644 2932
rect 1482 2892 1644 2898
rect 1992 2932 2154 2948
rect 1992 2898 2008 2932
rect 2042 2898 2154 2932
rect 1482 2882 1584 2892
rect 1992 2882 2154 2898
rect 3302 2932 3560 2948
rect 3302 2898 3318 2932
rect 3352 2898 3510 2932
rect 3544 2898 3560 2932
rect 3302 2882 3560 2898
rect 3912 2932 4170 2948
rect 3912 2898 3928 2932
rect 3962 2898 4120 2932
rect 4154 2898 4170 2932
rect 3912 2882 4170 2898
rect 5102 2932 5264 2948
rect 5102 2898 5118 2932
rect 5152 2898 5264 2932
rect 5102 2882 5264 2898
rect 5802 2932 5964 2948
rect 5802 2898 5818 2932
rect 5852 2898 5964 2932
rect 5802 2882 5964 2898
rect 1540 2428 1644 2438
rect 2054 2428 2154 2438
rect 1482 2422 1644 2428
rect 1482 2388 1594 2422
rect 1628 2388 1644 2422
rect 1482 2382 1644 2388
rect 1992 2422 2154 2428
rect 1992 2388 2104 2422
rect 2138 2388 2154 2422
rect 1992 2382 2154 2388
rect 1540 2372 1644 2382
rect 2054 2372 2154 2382
rect 3302 2422 3560 2438
rect 3302 2388 3414 2422
rect 3448 2388 3560 2422
rect 3302 2372 3560 2388
rect 3912 2422 4170 2438
rect 3912 2388 4024 2422
rect 4058 2388 4170 2422
rect 3912 2372 4170 2388
rect 5102 2422 5264 2438
rect 5102 2388 5214 2422
rect 5248 2388 5264 2422
rect 5102 2372 5264 2388
rect 5802 2422 5964 2438
rect 5802 2388 5914 2422
rect 5948 2388 5964 2422
rect 5802 2372 5964 2388
<< polycont >>
rect 1498 3736 1532 3770
rect 2008 3736 2042 3770
rect 3208 3736 3242 3770
rect 3400 3736 3434 3770
rect 3908 3736 3942 3770
rect 4100 3736 4134 3770
rect 4608 3736 4642 3770
rect 5118 3736 5152 3770
rect 5310 3736 5344 3770
rect 5818 3736 5852 3770
rect 6010 3736 6044 3770
rect 1594 3208 1628 3242
rect 2104 3208 2138 3242
rect 3304 3208 3338 3242
rect 3496 3208 3530 3242
rect 4004 3208 4038 3242
rect 4196 3208 4230 3242
rect 4704 3208 4738 3242
rect 5214 3208 5248 3242
rect 5406 3208 5440 3242
rect 5914 3208 5948 3242
rect 6106 3208 6140 3242
rect 1498 2898 1532 2932
rect 2008 2898 2042 2932
rect 3318 2898 3352 2932
rect 3510 2898 3544 2932
rect 3928 2898 3962 2932
rect 4120 2898 4154 2932
rect 5118 2898 5152 2932
rect 5818 2898 5852 2932
rect 1594 2388 1628 2422
rect 2104 2388 2138 2422
rect 3414 2388 3448 2422
rect 4024 2388 4058 2422
rect 5214 2388 5248 2422
rect 5914 2388 5948 2422
<< locali >>
rect 1780 3850 1870 3870
rect 1482 3736 1498 3770
rect 1532 3736 1644 3770
rect 1770 3630 1780 3760
rect 1860 3790 1870 3850
rect 3680 3780 3770 3870
rect 1992 3736 2008 3770
rect 2042 3736 2154 3770
rect 3192 3736 3208 3770
rect 3242 3736 3400 3770
rect 3434 3736 3546 3770
rect 1260 3240 1350 3530
rect 1770 3440 1860 3630
rect 3700 3540 3770 3780
rect 3892 3736 3908 3770
rect 3942 3736 4100 3770
rect 4134 3736 4246 3770
rect 1480 3242 1650 3250
rect 1260 3110 1360 3240
rect 1480 3208 1594 3242
rect 1628 3208 1650 3242
rect 1480 3200 1650 3208
rect 1780 3240 1860 3440
rect 1780 3110 1870 3240
rect 1992 3208 2104 3242
rect 2138 3208 2154 3242
rect 2290 3240 2370 3530
rect 2290 3110 2390 3240
rect 3192 3208 3304 3242
rect 3338 3208 3496 3242
rect 3530 3208 3546 3242
rect 3680 3110 3770 3540
rect 3892 3208 4004 3242
rect 4038 3208 4196 3242
rect 4230 3208 4246 3242
rect 4380 3110 4460 3870
rect 4592 3736 4608 3770
rect 4642 3736 4754 3770
rect 4592 3208 4704 3242
rect 4738 3208 4754 3242
rect 4890 3110 4970 3870
rect 5102 3736 5118 3770
rect 5152 3736 5310 3770
rect 5344 3736 5456 3770
rect 5102 3208 5214 3242
rect 5248 3208 5406 3242
rect 5440 3208 5456 3242
rect 5590 3110 5670 3870
rect 5802 3736 5818 3770
rect 5852 3736 6010 3770
rect 6044 3736 6156 3770
rect 5802 3208 5914 3242
rect 5948 3208 6106 3242
rect 6140 3208 6156 3242
rect 1482 2898 1498 2932
rect 1532 2898 1644 2932
rect 1770 2890 1870 3030
rect 1992 2898 2008 2932
rect 2042 2898 2154 2932
rect 3302 2898 3318 2932
rect 3352 2898 3510 2932
rect 3544 2898 3560 2932
rect 1770 2560 1860 2890
rect 1482 2388 1594 2422
rect 1628 2388 1644 2422
rect 1770 2310 1870 2560
rect 1992 2388 2104 2422
rect 2138 2388 2154 2422
rect 3302 2388 3414 2422
rect 3448 2388 3560 2422
rect 1340 2210 1750 2300
rect 1890 2260 3330 2300
rect 3530 2260 3580 2300
rect 3700 2290 3780 3030
rect 3912 2898 3928 2932
rect 3962 2898 4120 2932
rect 4154 2898 4170 2932
rect 5102 2898 5118 2932
rect 5152 2898 5264 2932
rect 5802 2898 5818 2932
rect 5852 2898 5964 2932
rect 3912 2388 4024 2422
rect 4058 2388 4170 2422
rect 5102 2388 5214 2422
rect 5248 2388 5264 2422
rect 5802 2388 5914 2422
rect 5948 2388 5964 2422
rect 1890 2210 3580 2260
rect 2250 2200 3580 2210
<< viali >>
rect 1498 3736 1532 3770
rect 1780 3630 1860 3850
rect 3960 3820 4160 3900
rect 2008 3736 2042 3770
rect 3208 3736 3242 3770
rect 3400 3736 3434 3770
rect 1250 3530 1360 3610
rect 2270 3530 2380 3610
rect 3640 3540 3700 3780
rect 3908 3736 3942 3770
rect 4100 3736 4134 3770
rect 1594 3208 1628 3242
rect 2104 3208 2138 3242
rect 3304 3208 3338 3242
rect 3496 3208 3530 3242
rect 4004 3208 4038 3242
rect 4196 3208 4230 3242
rect 4570 3820 4770 3900
rect 4608 3736 4642 3770
rect 4704 3208 4738 3242
rect 5180 3820 5380 3900
rect 5118 3736 5152 3770
rect 5310 3736 5344 3770
rect 5214 3208 5248 3242
rect 5406 3208 5440 3242
rect 5880 3820 6080 3900
rect 5818 3736 5852 3770
rect 6010 3736 6044 3770
rect 5914 3208 5948 3242
rect 6106 3208 6140 3242
rect 1498 2898 1532 2932
rect 2008 2898 2042 2932
rect 3318 2898 3352 2932
rect 3510 2898 3544 2932
rect 1594 2388 1628 2422
rect 2104 2388 2138 2422
rect 3414 2388 3448 2422
rect 1750 2210 1890 2310
rect 3330 2260 3530 2340
rect 3928 2898 3962 2932
rect 4120 2898 4154 2932
rect 5118 2898 5152 2932
rect 5818 2898 5852 2932
rect 4024 2388 4058 2422
rect 5214 2388 5248 2422
rect 5914 2388 5948 2422
rect 3940 2260 4140 2340
rect 4540 2260 4700 2340
rect 5090 2260 5290 2340
rect 5780 2260 5980 2340
rect 1740 1460 1910 1530
<< metal1 >>
rect 3948 3900 4172 3906
rect 1774 3860 1866 3862
rect 1482 3770 1644 3776
rect 1482 3736 1498 3770
rect 1532 3736 1644 3770
rect 1740 3740 1750 3860
rect 1890 3740 1900 3860
rect 2490 3820 3790 3870
rect 1992 3770 2154 3776
rect 1482 3730 1644 3736
rect 1238 3610 1372 3616
rect 1238 3530 1250 3610
rect 1360 3530 1372 3610
rect 1238 3524 1372 3530
rect 1430 3512 1440 3688
rect 1494 3512 1504 3688
rect 1070 3430 1320 3480
rect 1540 3466 1590 3730
rect 1622 3512 1632 3688
rect 1686 3512 1696 3688
rect 1774 3630 1780 3740
rect 1860 3630 1866 3740
rect 1992 3736 2008 3770
rect 2042 3736 2154 3770
rect 1992 3730 2154 3736
rect 1774 3618 1866 3630
rect 1940 3512 1950 3688
rect 2004 3512 2014 3688
rect 2050 3466 2100 3730
rect 2132 3512 2142 3688
rect 2196 3512 2206 3688
rect 2258 3610 2392 3616
rect 2258 3530 2270 3610
rect 2380 3530 2392 3610
rect 2258 3524 2392 3530
rect 2490 3480 2550 3820
rect 3634 3780 3706 3792
rect 3740 3780 3790 3820
rect 3948 3820 3960 3900
rect 4160 3820 4172 3900
rect 3948 3814 4172 3820
rect 4558 3900 4782 3906
rect 4558 3820 4570 3900
rect 4770 3820 4782 3900
rect 4558 3814 4782 3820
rect 5168 3900 5392 3906
rect 5168 3820 5180 3900
rect 5380 3820 5392 3900
rect 5168 3814 5392 3820
rect 5868 3900 6092 3906
rect 5868 3820 5880 3900
rect 6080 3820 6092 3900
rect 5868 3814 6092 3820
rect 3040 3770 3550 3780
rect 3040 3736 3208 3770
rect 3242 3736 3400 3770
rect 3434 3736 3550 3770
rect 3040 3730 3550 3736
rect 910 3290 920 3390
rect 1080 3290 1090 3390
rect 1120 3290 1130 3390
rect 1230 3290 1240 3390
rect 1270 3250 1320 3430
rect 1526 3290 1536 3466
rect 1590 3290 1600 3466
rect 2036 3290 2046 3466
rect 2100 3290 2110 3466
rect 2310 3430 2570 3480
rect 1540 3250 1590 3290
rect 2050 3250 2100 3290
rect 2310 3250 2360 3430
rect 2390 3290 2400 3390
rect 2500 3290 2510 3390
rect 2540 3290 2550 3390
rect 2710 3290 2720 3390
rect 3040 3250 3090 3730
rect 3140 3514 3150 3690
rect 3204 3514 3214 3690
rect 3332 3514 3342 3690
rect 3396 3514 3406 3690
rect 3524 3514 3534 3690
rect 3588 3514 3598 3690
rect 3630 3540 3640 3780
rect 3700 3540 3710 3780
rect 3740 3770 4250 3780
rect 3740 3736 3908 3770
rect 3942 3736 4100 3770
rect 4134 3736 4250 3770
rect 3740 3730 4250 3736
rect 4440 3770 4760 3780
rect 4440 3736 4608 3770
rect 4642 3736 4760 3770
rect 4440 3730 4760 3736
rect 4950 3770 5460 3780
rect 4950 3736 5118 3770
rect 5152 3736 5310 3770
rect 5344 3736 5460 3770
rect 4950 3730 5460 3736
rect 5650 3770 6160 3780
rect 5650 3736 5818 3770
rect 5852 3736 6010 3770
rect 6044 3736 6160 3770
rect 5650 3730 6160 3736
rect 3634 3528 3706 3540
rect 3236 3288 3246 3464
rect 3300 3288 3310 3464
rect 3428 3288 3438 3464
rect 3492 3288 3502 3464
rect 3740 3250 3790 3730
rect 3840 3514 3850 3690
rect 3904 3514 3914 3690
rect 4032 3514 4042 3690
rect 4096 3514 4106 3690
rect 4224 3514 4234 3690
rect 4288 3514 4298 3690
rect 3936 3288 3946 3464
rect 4000 3288 4010 3464
rect 4128 3288 4138 3464
rect 4192 3288 4202 3464
rect 4440 3250 4500 3730
rect 4540 3514 4550 3690
rect 4604 3514 4614 3690
rect 4732 3514 4742 3690
rect 4796 3514 4806 3690
rect 4636 3288 4646 3464
rect 4700 3288 4710 3464
rect 4950 3250 5000 3730
rect 5050 3514 5060 3690
rect 5114 3514 5124 3690
rect 5242 3514 5252 3690
rect 5306 3514 5316 3690
rect 5434 3514 5444 3690
rect 5498 3514 5508 3690
rect 5146 3288 5156 3464
rect 5210 3288 5220 3464
rect 5338 3288 5348 3464
rect 5402 3288 5412 3464
rect 5650 3250 5700 3730
rect 5750 3514 5760 3690
rect 5814 3514 5824 3690
rect 5942 3514 5952 3690
rect 6006 3514 6016 3690
rect 6134 3514 6144 3690
rect 6198 3514 6208 3690
rect 5846 3288 5856 3464
rect 5910 3288 5920 3464
rect 6038 3286 6048 3462
rect 6102 3286 6112 3462
rect 1070 3200 1460 3250
rect 1450 3160 1460 3200
rect 1670 3160 1680 3250
rect 1960 3160 1970 3250
rect 2180 3200 2570 3250
rect 3040 3242 3550 3250
rect 3040 3208 3304 3242
rect 3338 3208 3496 3242
rect 3530 3208 3550 3242
rect 3040 3200 3550 3208
rect 3740 3242 4250 3250
rect 3740 3208 4004 3242
rect 4038 3208 4196 3242
rect 4230 3208 4250 3242
rect 3740 3200 4250 3208
rect 4440 3242 4760 3250
rect 4440 3208 4704 3242
rect 4738 3208 4760 3242
rect 4440 3200 4760 3208
rect 4950 3242 5460 3250
rect 4950 3208 5214 3242
rect 5248 3208 5406 3242
rect 5440 3208 5460 3242
rect 4950 3200 5460 3208
rect 5650 3242 6160 3250
rect 5650 3208 5914 3242
rect 5948 3208 6106 3242
rect 6140 3208 6160 3242
rect 5650 3200 6160 3208
rect 2180 3160 2190 3200
rect 1620 3120 1680 3160
rect 3040 3120 3090 3200
rect 4440 3150 4500 3200
rect 4950 3150 5000 3200
rect 5650 3150 5700 3200
rect 1620 3070 3090 3120
rect 1330 2932 1650 2950
rect 1330 2898 1498 2932
rect 1532 2898 1650 2932
rect 1330 2890 1650 2898
rect 1990 2932 2310 2950
rect 1990 2898 2008 2932
rect 2042 2898 2310 2932
rect 1990 2890 2310 2898
rect 3290 2920 3300 3010
rect 3560 2940 3570 3010
rect 4430 3000 4440 3150
rect 4510 3000 4520 3150
rect 4940 3000 4950 3150
rect 5010 3000 5020 3150
rect 5640 3000 5650 3150
rect 5710 3000 5720 3150
rect 4440 2940 4500 3000
rect 4950 2940 5000 3000
rect 5650 2940 5700 3000
rect 3560 2932 4180 2940
rect 3560 2920 3928 2932
rect 3290 2898 3318 2920
rect 3352 2898 3510 2920
rect 3544 2898 3928 2920
rect 3962 2898 4120 2932
rect 4154 2898 4180 2932
rect 3290 2890 4180 2898
rect 4440 2890 4660 2940
rect 4950 2932 5270 2940
rect 4950 2898 5118 2932
rect 5152 2898 5270 2932
rect 4950 2890 5270 2898
rect 5650 2932 5970 2940
rect 5650 2898 5818 2932
rect 5852 2898 5970 2932
rect 5650 2890 5970 2898
rect 1330 2430 1390 2890
rect 1526 2684 1536 2860
rect 1590 2684 1600 2860
rect 2036 2684 2046 2860
rect 2100 2684 2110 2860
rect 1430 2460 1440 2636
rect 1494 2460 1504 2636
rect 1622 2460 1632 2636
rect 1686 2460 1696 2636
rect 1940 2460 1950 2636
rect 2004 2460 2014 2636
rect 2132 2460 2142 2636
rect 2196 2460 2206 2636
rect 2250 2430 2310 2890
rect 3346 2684 3356 2860
rect 3410 2684 3420 2860
rect 3538 2684 3548 2860
rect 3602 2684 3612 2860
rect 3250 2460 3260 2636
rect 3314 2460 3324 2636
rect 3442 2460 3452 2636
rect 3506 2460 3516 2636
rect 3710 2430 3760 2890
rect 3956 2684 3966 2860
rect 4020 2684 4030 2860
rect 4148 2684 4158 2860
rect 4212 2684 4222 2860
rect 3860 2460 3870 2636
rect 3924 2460 3934 2636
rect 4052 2460 4062 2636
rect 4116 2460 4126 2636
rect 4440 2430 4500 2890
rect 4628 2684 4638 2860
rect 4692 2684 4702 2860
rect 4540 2460 4550 2636
rect 4604 2460 4614 2636
rect 4950 2430 5000 2890
rect 5146 2684 5156 2860
rect 5210 2684 5220 2860
rect 5050 2460 5060 2636
rect 5114 2460 5124 2636
rect 5242 2460 5252 2636
rect 5306 2460 5316 2636
rect 5650 2430 5700 2890
rect 5846 2684 5856 2860
rect 5910 2684 5920 2860
rect 5750 2460 5760 2636
rect 5814 2460 5824 2636
rect 5942 2460 5952 2636
rect 6006 2460 6016 2636
rect 1330 2422 1650 2430
rect 1330 2388 1594 2422
rect 1628 2388 1650 2422
rect 1330 2370 1650 2388
rect 1990 2422 2310 2430
rect 1990 2388 2104 2422
rect 2138 2388 2310 2422
rect 1990 2370 2310 2388
rect 3290 2422 4180 2430
rect 3290 2388 3414 2422
rect 3448 2388 4024 2422
rect 4058 2388 4180 2422
rect 3290 2380 4180 2388
rect 4440 2380 4660 2430
rect 4950 2422 5270 2430
rect 4950 2388 5214 2422
rect 5248 2388 5270 2422
rect 4950 2380 5270 2388
rect 5650 2422 5970 2430
rect 5650 2388 5914 2422
rect 5948 2388 5970 2422
rect 5650 2380 5970 2388
rect 3318 2340 3542 2346
rect 1738 2310 1902 2316
rect 3318 2310 3330 2340
rect 1738 2210 1750 2310
rect 1890 2260 3330 2310
rect 3530 2260 3542 2340
rect 1890 2254 3542 2260
rect 3928 2340 4152 2346
rect 3928 2260 3940 2340
rect 4140 2260 4152 2340
rect 3928 2254 4152 2260
rect 4528 2340 4712 2346
rect 4528 2260 4540 2340
rect 4700 2260 4712 2340
rect 4528 2254 4712 2260
rect 5078 2340 5302 2346
rect 5078 2260 5090 2340
rect 5290 2260 5302 2340
rect 5078 2254 5302 2260
rect 5768 2340 5992 2346
rect 5768 2260 5780 2340
rect 5980 2260 5992 2340
rect 5768 2254 5992 2260
rect 1890 2210 3530 2254
rect 1738 2204 1902 2210
rect 1070 2050 1190 2130
rect 1230 2080 3310 2130
rect 1050 1874 1060 2050
rect 1114 1874 1190 2050
rect 1070 1826 1190 1874
rect 1280 2050 1370 2080
rect 3340 2050 3480 2130
rect 1280 1874 1296 2050
rect 1350 1874 1370 2050
rect 1522 1874 1532 2050
rect 1586 1874 1596 2050
rect 1758 1874 1768 2050
rect 1822 1874 1832 2050
rect 1994 1874 2004 2050
rect 2058 1874 2068 2050
rect 2230 1874 2240 2050
rect 2294 1874 2304 2050
rect 2466 1874 2476 2050
rect 2530 1874 2540 2050
rect 2702 1874 2712 2050
rect 2766 1874 2776 2050
rect 2938 1874 2948 2050
rect 3002 1874 3012 2050
rect 3174 1874 3184 2050
rect 3238 1874 3248 2050
rect 3340 1874 3420 2050
rect 3474 1874 3484 2050
rect 1070 1650 1178 1826
rect 1232 1650 1242 1826
rect 1070 1570 1190 1650
rect 1280 1620 1370 1874
rect 3340 1826 3480 1874
rect 1404 1650 1414 1826
rect 1468 1650 1478 1826
rect 1640 1650 1650 1826
rect 1704 1650 1714 1826
rect 1876 1650 1886 1826
rect 1940 1650 1950 1826
rect 2112 1650 2122 1826
rect 2176 1650 2186 1826
rect 2348 1650 2358 1826
rect 2412 1650 2422 1826
rect 2584 1650 2594 1826
rect 2648 1650 2658 1826
rect 2820 1650 2830 1826
rect 2884 1650 2894 1826
rect 3056 1650 3066 1826
rect 3120 1650 3130 1826
rect 3292 1650 3302 1826
rect 3356 1650 3480 1826
rect 1230 1570 3310 1620
rect 3340 1570 3480 1650
rect 1728 1530 1922 1536
rect 1728 1460 1740 1530
rect 1910 1460 1922 1530
rect 1728 1454 1922 1460
<< via1 >>
rect 1750 3850 1890 3860
rect 1750 3740 1780 3850
rect 1780 3740 1860 3850
rect 1860 3740 1890 3850
rect 1250 3530 1360 3610
rect 1440 3512 1494 3688
rect 1632 3512 1686 3688
rect 1950 3512 2004 3688
rect 2142 3512 2196 3688
rect 2270 3530 2380 3610
rect 3960 3820 4160 3900
rect 4570 3820 4770 3900
rect 5180 3820 5380 3900
rect 5880 3820 6080 3900
rect 920 3290 1080 3390
rect 1130 3290 1230 3390
rect 1536 3290 1590 3466
rect 2046 3290 2100 3466
rect 2400 3290 2500 3390
rect 2550 3290 2710 3390
rect 3150 3514 3204 3690
rect 3342 3514 3396 3690
rect 3534 3514 3588 3690
rect 3640 3540 3700 3780
rect 3246 3288 3300 3464
rect 3438 3288 3492 3464
rect 3850 3514 3904 3690
rect 4042 3514 4096 3690
rect 4234 3514 4288 3690
rect 3946 3288 4000 3464
rect 4138 3288 4192 3464
rect 4550 3514 4604 3690
rect 4742 3514 4796 3690
rect 4646 3288 4700 3464
rect 5060 3514 5114 3690
rect 5252 3514 5306 3690
rect 5444 3514 5498 3690
rect 5156 3288 5210 3464
rect 5348 3288 5402 3464
rect 5760 3514 5814 3690
rect 5952 3514 6006 3690
rect 6144 3514 6198 3690
rect 5856 3288 5910 3464
rect 6048 3286 6102 3462
rect 1460 3242 1670 3250
rect 1460 3208 1594 3242
rect 1594 3208 1628 3242
rect 1628 3208 1670 3242
rect 1460 3160 1670 3208
rect 1970 3242 2180 3250
rect 1970 3208 2104 3242
rect 2104 3208 2138 3242
rect 2138 3208 2180 3242
rect 1970 3160 2180 3208
rect 3300 2932 3560 3010
rect 4440 3000 4510 3150
rect 4950 3000 5010 3150
rect 5650 3000 5710 3150
rect 3300 2920 3318 2932
rect 3318 2920 3352 2932
rect 3352 2920 3510 2932
rect 3510 2920 3544 2932
rect 3544 2920 3560 2932
rect 1536 2684 1590 2860
rect 2046 2684 2100 2860
rect 1440 2460 1494 2636
rect 1632 2460 1686 2636
rect 1950 2460 2004 2636
rect 2142 2460 2196 2636
rect 3356 2684 3410 2860
rect 3548 2684 3602 2860
rect 3260 2460 3314 2636
rect 3452 2460 3506 2636
rect 3966 2684 4020 2860
rect 4158 2684 4212 2860
rect 3870 2460 3924 2636
rect 4062 2460 4116 2636
rect 4638 2684 4692 2860
rect 4550 2460 4604 2636
rect 5156 2684 5210 2860
rect 5060 2460 5114 2636
rect 5252 2460 5306 2636
rect 5856 2684 5910 2860
rect 5760 2460 5814 2636
rect 5952 2460 6006 2636
rect 3330 2260 3530 2340
rect 3940 2260 4140 2340
rect 4540 2260 4700 2340
rect 5090 2260 5290 2340
rect 5780 2260 5980 2340
rect 1060 1874 1114 2050
rect 1296 1874 1350 2050
rect 1532 1874 1586 2050
rect 1768 1874 1822 2050
rect 2004 1874 2058 2050
rect 2240 1874 2294 2050
rect 2476 1874 2530 2050
rect 2712 1874 2766 2050
rect 2948 1874 3002 2050
rect 3184 1874 3238 2050
rect 3420 1874 3474 2050
rect 1178 1650 1232 1826
rect 1414 1650 1468 1826
rect 1650 1650 1704 1826
rect 1886 1650 1940 1826
rect 2122 1650 2176 1826
rect 2358 1650 2412 1826
rect 2594 1650 2648 1826
rect 2830 1650 2884 1826
rect 3066 1650 3120 1826
rect 3302 1650 3356 1826
rect 1740 1460 1910 1530
<< metal2 >>
rect 920 3900 6340 3910
rect 920 3860 3960 3900
rect 920 3740 1750 3860
rect 1890 3820 3960 3860
rect 4160 3820 4570 3900
rect 4770 3820 5180 3900
rect 5380 3820 5880 3900
rect 6080 3820 6340 3900
rect 1890 3780 6340 3820
rect 1890 3740 3640 3780
rect 920 3690 3640 3740
rect 920 3688 1710 3690
rect 920 3610 1440 3688
rect 920 3530 1250 3610
rect 1360 3530 1440 3610
rect 920 3390 1080 3530
rect 1250 3520 1360 3530
rect 1494 3530 1632 3688
rect 1440 3502 1494 3512
rect 1686 3530 1710 3688
rect 1930 3688 3150 3690
rect 1930 3530 1950 3688
rect 1632 3502 1686 3512
rect 2004 3530 2142 3688
rect 1950 3502 2004 3512
rect 2196 3610 3150 3688
rect 2196 3530 2270 3610
rect 2380 3560 3150 3610
rect 2380 3530 2710 3560
rect 2270 3520 2380 3530
rect 2142 3502 2196 3512
rect 1536 3466 1590 3476
rect 920 3280 1080 3290
rect 1130 3400 1230 3410
rect 1130 3270 1230 3280
rect 1460 3290 1536 3440
rect 2046 3466 2100 3476
rect 1590 3290 1670 3440
rect 1460 3250 1670 3290
rect 1460 3130 1670 3160
rect 1460 3010 1560 3130
rect 1460 2860 1670 3010
rect 1460 2710 1536 2860
rect 1590 2710 1670 2860
rect 1970 3320 2046 3440
rect 2100 3290 2180 3440
rect 2080 3250 2180 3290
rect 2400 3400 2500 3410
rect 2550 3390 2710 3530
rect 3204 3560 3342 3690
rect 3150 3504 3204 3514
rect 3396 3560 3534 3690
rect 3342 3504 3396 3514
rect 3588 3560 3640 3690
rect 3700 3690 6340 3780
rect 3700 3560 3850 3690
rect 3640 3530 3700 3540
rect 3534 3504 3588 3514
rect 3904 3560 4042 3690
rect 3850 3504 3904 3514
rect 4096 3560 4234 3690
rect 4042 3504 4096 3514
rect 4288 3560 4550 3690
rect 4234 3504 4288 3514
rect 4604 3560 4742 3690
rect 4550 3504 4604 3514
rect 4796 3560 5060 3690
rect 4742 3504 4796 3514
rect 5114 3560 5252 3690
rect 5060 3504 5114 3514
rect 5306 3560 5444 3690
rect 5252 3504 5306 3514
rect 5498 3560 5760 3690
rect 5444 3504 5498 3514
rect 5814 3560 5952 3690
rect 5760 3504 5814 3514
rect 6006 3560 6144 3690
rect 5952 3504 6006 3514
rect 6198 3560 6340 3690
rect 6144 3504 6198 3514
rect 3246 3464 3300 3474
rect 2550 3280 2710 3290
rect 3190 3288 3246 3410
rect 3438 3464 3492 3474
rect 3300 3288 3438 3410
rect 3946 3464 4000 3474
rect 3492 3288 3570 3410
rect 2400 3270 2500 3280
rect 3190 3250 3570 3288
rect 1970 2860 2180 3160
rect 1970 2710 2046 2860
rect 1536 2674 1590 2684
rect 2100 2710 2180 2860
rect 3270 3010 3570 3250
rect 3270 2920 3300 3010
rect 3560 2920 3570 3010
rect 3270 2900 3570 2920
rect 3920 3288 3946 3410
rect 4138 3464 4192 3474
rect 4000 3288 4138 3410
rect 4646 3464 4700 3474
rect 4192 3288 4220 3410
rect 3920 3110 4220 3288
rect 4620 3288 4646 3430
rect 5156 3464 5210 3474
rect 4700 3288 4730 3430
rect 4440 3150 4510 3160
rect 3920 3050 4440 3110
rect 3270 2860 3650 2900
rect 3270 2740 3356 2860
rect 2046 2674 2100 2684
rect 3410 2740 3548 2860
rect 3356 2674 3410 2684
rect 3602 2740 3650 2860
rect 3920 2860 4220 3050
rect 4440 2990 4510 3000
rect 4620 3110 4730 3288
rect 5130 3288 5156 3440
rect 5348 3464 5402 3474
rect 5210 3288 5348 3440
rect 5856 3464 5910 3474
rect 5402 3288 5420 3440
rect 5130 3270 5420 3288
rect 5830 3288 5856 3440
rect 6048 3462 6102 3472
rect 5910 3288 6048 3440
rect 5830 3286 6048 3288
rect 6102 3286 6120 3440
rect 5830 3270 6120 3286
rect 4950 3150 5010 3160
rect 4620 3050 4950 3110
rect 3920 2740 3966 2860
rect 3548 2674 3602 2684
rect 4020 2740 4158 2860
rect 3966 2674 4020 2684
rect 4212 2740 4220 2860
rect 4620 2860 4730 3050
rect 4950 2990 5010 3000
rect 5130 3110 5240 3270
rect 5650 3150 5710 3160
rect 5130 3050 5650 3110
rect 4620 2720 4638 2860
rect 4158 2674 4212 2684
rect 4692 2720 4730 2860
rect 5130 2860 5240 3050
rect 5650 2990 5710 3000
rect 5130 2730 5156 2860
rect 4638 2674 4692 2684
rect 5210 2730 5240 2860
rect 5830 2860 5940 3270
rect 5830 2730 5856 2860
rect 5156 2674 5210 2684
rect 5910 2730 5940 2860
rect 5856 2674 5910 2684
rect 1440 2636 1494 2646
rect 1430 2460 1440 2610
rect 1632 2636 1686 2646
rect 1494 2460 1632 2610
rect 1950 2636 2004 2646
rect 1686 2460 1950 2610
rect 2142 2636 2196 2646
rect 2004 2460 2142 2610
rect 3260 2636 3314 2646
rect 2196 2460 2730 2610
rect 1430 2340 2730 2460
rect 3220 2460 3260 2590
rect 3452 2636 3506 2646
rect 3314 2460 3452 2590
rect 3870 2636 3924 2646
rect 3506 2460 3870 2590
rect 4062 2636 4116 2646
rect 3924 2460 4062 2590
rect 4550 2636 4604 2646
rect 4116 2460 4550 2590
rect 5060 2636 5114 2646
rect 4604 2460 5060 2590
rect 5252 2636 5306 2646
rect 5114 2460 5252 2590
rect 5760 2636 5814 2646
rect 5306 2460 5760 2590
rect 5952 2636 6006 2646
rect 5814 2460 5952 2590
rect 6006 2460 6050 2590
rect 3220 2410 6050 2460
rect 3310 2340 6050 2410
rect 1430 2250 3240 2340
rect 1050 2050 1120 2060
rect 1050 1874 1060 2050
rect 1114 1874 1120 2050
rect 1250 2050 1400 2160
rect 1250 1920 1296 2050
rect 1050 1780 1120 1874
rect 1350 1920 1400 2050
rect 1510 2050 3240 2250
rect 1510 1920 1532 2050
rect 1296 1864 1350 1874
rect 1586 1920 1768 2050
rect 1532 1864 1586 1874
rect 1822 1920 2004 2050
rect 1768 1864 1822 1874
rect 2058 1920 2240 2050
rect 2004 1864 2058 1874
rect 2294 1920 2476 2050
rect 2240 1864 2294 1874
rect 2530 1920 2712 2050
rect 2476 1864 2530 1874
rect 2766 1920 2948 2050
rect 2712 1864 2766 1874
rect 3002 1920 3184 2050
rect 2948 1864 3002 1874
rect 3238 1920 3240 2050
rect 3310 2260 3330 2340
rect 3530 2260 3940 2340
rect 4140 2260 4540 2340
rect 4700 2260 5090 2340
rect 5290 2260 5780 2340
rect 5980 2260 6050 2340
rect 3310 2250 6050 2260
rect 3310 2050 3640 2250
rect 3184 1864 3238 1874
rect 3310 1874 3420 2050
rect 3474 1874 3640 2050
rect 1178 1826 1232 1836
rect 1050 1650 1178 1780
rect 1414 1826 1468 1836
rect 1232 1650 1414 1780
rect 1650 1826 1704 1836
rect 1468 1650 1650 1780
rect 1886 1826 1940 1836
rect 1704 1650 1886 1780
rect 2122 1826 2176 1836
rect 1940 1650 2122 1780
rect 2358 1826 2412 1836
rect 2176 1650 2358 1780
rect 2594 1826 2648 1836
rect 2412 1650 2594 1780
rect 2830 1826 2884 1836
rect 2648 1650 2830 1780
rect 3066 1826 3120 1836
rect 3310 1830 3640 1874
rect 2884 1650 3066 1780
rect 3290 1826 3640 1830
rect 3290 1780 3302 1826
rect 3120 1650 3302 1780
rect 3356 1650 3640 1826
rect 1050 1530 3640 1650
rect 1050 1480 1740 1530
rect 1910 1480 3640 1530
rect 1740 1450 1910 1460
<< via2 >>
rect 1130 3390 1230 3400
rect 1130 3290 1230 3390
rect 1130 3280 1230 3290
rect 1560 3010 1670 3130
rect 1970 3290 2046 3320
rect 2046 3290 2080 3320
rect 1970 3250 2080 3290
rect 2400 3390 2500 3400
rect 2400 3290 2500 3390
rect 2400 3280 2500 3290
rect 1970 3200 2080 3250
<< metal3 >>
rect 1120 3400 1240 3405
rect 2390 3400 2510 3405
rect 1120 3280 1130 3400
rect 1230 3320 1370 3400
rect 1960 3320 2090 3325
rect 1230 3280 1970 3320
rect 1120 3275 1970 3280
rect 1220 3200 1970 3275
rect 2080 3200 2090 3320
rect 2390 3280 2400 3400
rect 2500 3280 2510 3400
rect 2390 3275 2510 3280
rect 1960 3195 2090 3200
rect 1550 3130 1680 3135
rect 2400 3130 2500 3275
rect 1550 3010 1560 3130
rect 1670 3010 2500 3130
rect 1550 3005 1680 3010
use sky130_fd_pr__nfet_01v8_GV8PGY  sky130_fd_pr__nfet_01v8_GV8PGY_0
timestamp 1654768133
transform 1 0 3431 0 1 2660
box -311 -410 311 410
use sky130_fd_pr__nfet_01v8_GV8PGY  sky130_fd_pr__nfet_01v8_GV8PGY_1
timestamp 1654768133
transform 1 0 4041 0 1 2660
box -311 -410 311 410
use sky130_fd_pr__nfet_01v8_PL8DH5  sky130_fd_pr__nfet_01v8_PL8DH5_0
timestamp 1654768133
transform 1 0 2267 0 1 1850
box -1347 -410 1347 410
use sky130_fd_pr__nfet_01v8_YT8PGU  sky130_fd_pr__nfet_01v8_YT8PGU_0
timestamp 1654768133
transform 1 0 4621 0 1 2660
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_lvt_LH2JGW  sky130_fd_pr__nfet_01v8_lvt_LH2JGW_0
timestamp 1654768133
transform 1 0 1563 0 1 2660
box -263 -410 263 410
use sky130_fd_pr__nfet_01v8_lvt_LH2JGW  sky130_fd_pr__nfet_01v8_lvt_LH2JGW_1
timestamp 1654768133
transform 1 0 2073 0 1 2660
box -263 -410 263 410
use sky130_fd_pr__nfet_01v8_lvt_LH2JGW  sky130_fd_pr__nfet_01v8_lvt_LH2JGW_2
timestamp 1654768133
transform 1 0 5883 0 1 2660
box -263 -410 263 410
use sky130_fd_pr__nfet_01v8_lvt_LH2JGW  sky130_fd_pr__nfet_01v8_lvt_LH2JGW_3
timestamp 1654768133
transform 1 0 5183 0 1 2660
box -263 -410 263 410
use sky130_fd_pr__pfet_01v8_U47ZGH  sky130_fd_pr__pfet_01v8_U47ZGH_0
timestamp 1654768133
transform 1 0 3369 0 1 3489
box -359 -419 359 419
use sky130_fd_pr__pfet_01v8_U47ZGH  sky130_fd_pr__pfet_01v8_U47ZGH_1
timestamp 1654768133
transform 1 0 4069 0 1 3489
box -359 -419 359 419
use sky130_fd_pr__pfet_01v8_U47ZGH  sky130_fd_pr__pfet_01v8_U47ZGH_2
timestamp 1654768133
transform 1 0 5279 0 1 3489
box -359 -419 359 419
use sky130_fd_pr__pfet_01v8_U47ZGH  sky130_fd_pr__pfet_01v8_U47ZGH_3
timestamp 1654768133
transform 1 0 5979 0 1 3489
box -359 -419 359 419
use sky130_fd_pr__pfet_01v8_X4XKHL  sky130_fd_pr__pfet_01v8_X4XKHL_0
timestamp 1654768133
transform 1 0 1563 0 1 3489
box -263 -419 263 419
use sky130_fd_pr__pfet_01v8_X4XKHL  sky130_fd_pr__pfet_01v8_X4XKHL_1
timestamp 1654768133
transform 1 0 2073 0 1 3489
box -263 -419 263 419
use sky130_fd_pr__pfet_01v8_X4XKHL  sky130_fd_pr__pfet_01v8_X4XKHL_2
timestamp 1654768133
transform 1 0 4673 0 1 3489
box -263 -419 263 419
use sky130_fd_pr__pfet_01v8_XJ7GBL  sky130_fd_pr__pfet_01v8_XJ7GBL_0
timestamp 1654768133
transform 1 0 1101 0 1 3339
box -211 -269 211 269
use sky130_fd_pr__pfet_01v8_XJ7GBL  sky130_fd_pr__pfet_01v8_XJ7GBL_1
timestamp 1654768133
transform 1 0 2531 0 1 3339
box -211 -269 211 269
<< labels >>
rlabel metal2 5850 3020 5930 3130 1 Out
rlabel metal2 1250 1920 1400 2160 1 I_Bias
rlabel metal1 1330 2580 1390 2780 1 In_n
rlabel metal1 2250 2580 2310 2780 1 In_p
rlabel metal2 2650 3660 2850 3760 1 VP
rlabel metal2 5550 3050 5610 3110 1 VM13D
rlabel metal2 4850 3050 4910 3110 1 VM17D
rlabel metal2 4340 3050 4400 3110 1 VM12D
rlabel metal2 3370 3050 3430 3110 1 VM11D
rlabel metal2 1530 2980 1590 3040 1 VM1D
rlabel metal2 2050 2980 2110 3040 1 VM6D
rlabel metal2 1790 2220 1850 2280 1 VM4D
rlabel metal2 3458 2114 3576 2222 1 VN
<< end >>
