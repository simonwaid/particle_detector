magic
tech sky130A
magscale 1 2
timestamp 1654695234
<< nwell >>
rect 2940 6920 6680 7160
rect 660 6100 6340 6260
rect 660 5830 1230 6100
rect 1250 5830 6340 6100
rect 660 5820 6340 5830
rect 2920 5090 6640 5330
rect 650 3990 6320 4430
<< pwell >>
rect 2980 6390 6300 6610
rect 2980 6380 6250 6390
rect 2980 6310 6310 6380
rect 6220 6300 6310 6310
rect 660 5410 6310 5740
rect 16060 5170 20880 5240
rect 20790 5120 20880 5170
rect 17420 4960 17550 5010
rect 2960 4560 6280 4780
rect 2960 4550 6230 4560
rect 2960 4480 6290 4550
rect 6200 4470 6290 4480
rect 650 3900 6320 3910
rect 650 3730 800 3900
rect 880 3730 6320 3900
rect 650 3580 6320 3730
<< psubdiff >>
rect 3010 6360 6280 6370
rect 3010 6320 3040 6360
rect 6250 6320 6280 6360
rect 3010 6310 6280 6320
rect 660 5430 700 5500
rect 6250 5430 6310 5500
rect 660 5410 6310 5430
rect 2990 4530 6260 4540
rect 2990 4490 3020 4530
rect 6230 4490 6260 4530
rect 2990 4480 6260 4490
rect 650 3610 690 3670
rect 6270 3610 6320 3670
rect 650 3580 6320 3610
<< nsubdiff >>
rect 2980 7080 6340 7120
rect 2980 7040 3040 7080
rect 6280 7040 6340 7080
rect 2980 7010 6340 7040
rect 700 6190 1200 6210
rect 700 6150 730 6190
rect 1170 6150 1200 6190
rect 700 6140 1200 6150
rect 1270 6200 6270 6220
rect 1270 6160 1310 6200
rect 6240 6160 6270 6200
rect 1270 6140 6270 6160
rect 2960 5250 6320 5290
rect 2960 5210 3020 5250
rect 6260 5210 6320 5250
rect 2960 5180 6320 5210
rect 690 4360 1190 4380
rect 690 4320 720 4360
rect 1160 4320 1190 4360
rect 690 4310 1190 4320
rect 1250 4370 6250 4390
rect 1250 4330 1290 4370
rect 6220 4330 6250 4370
rect 1250 4310 6250 4330
<< psubdiffcont >>
rect 3040 6320 6250 6360
rect 700 5430 6250 5500
rect 3020 4490 6230 4530
rect 690 3610 6270 3670
<< nsubdiffcont >>
rect 3040 7040 6280 7080
rect 730 6150 1170 6190
rect 1310 6160 6240 6200
rect 3020 5210 6260 5250
rect 720 4320 1160 4360
rect 1290 4330 6220 4370
<< locali >>
rect 3440 11840 3530 20040
rect 5170 11840 5270 20040
rect 6910 11840 7010 20040
rect 10390 11840 10490 20040
rect 12130 11840 12230 20040
rect 13870 11840 13970 20040
rect 15610 11840 15710 20040
rect 17350 11840 17450 20040
rect 3440 10270 3530 11610
rect 3340 10250 3530 10270
rect 5170 10260 5270 11610
rect 6910 10260 7010 11610
rect 10390 10260 10490 11610
rect 12130 10260 12230 11610
rect 13870 10260 13970 11610
rect 15610 10260 15710 11610
rect 17350 10630 17450 11610
rect 17350 10260 17450 10300
rect 19090 10260 19190 11610
rect 3340 7530 3510 10250
rect 6650 7120 13560 7540
rect 2980 7080 6310 7100
rect 2980 7040 3040 7080
rect 6280 7040 6310 7080
rect 2980 7030 6310 7040
rect 3010 6360 6310 6380
rect 3010 6320 3040 6360
rect 6250 6320 6310 6360
rect 3010 6300 6310 6320
rect 700 6190 1200 6210
rect 700 6150 730 6190
rect 1170 6150 1200 6190
rect 700 6140 1200 6150
rect 1270 6200 6270 6220
rect 1270 6160 1310 6200
rect 6240 6160 6270 6200
rect 1270 6140 6270 6160
rect 660 5430 700 5500
rect 6250 5430 6310 5500
rect 660 5410 6310 5430
rect 2960 5250 6290 5270
rect 2960 5210 3020 5250
rect 6260 5210 6290 5250
rect 2960 5200 6290 5210
rect 2990 4530 6290 4550
rect 2990 4490 3020 4530
rect 6230 4490 6290 4530
rect 2990 4470 6290 4490
rect 690 4360 1190 4380
rect 690 4320 720 4360
rect 1160 4320 1190 4360
rect 690 4310 1190 4320
rect 1250 4370 6250 4390
rect 1250 4330 1290 4370
rect 6220 4330 6250 4370
rect 1250 4310 6250 4330
rect 650 3610 690 3670
rect 6270 3610 6320 3670
rect 13080 3650 13680 4230
rect 14300 3650 14400 6740
rect 15000 3650 15300 6760
rect 15900 3650 16000 6780
rect 19100 3760 19180 5100
rect 17350 3650 20840 3760
rect 13080 3640 20840 3650
rect 650 3580 6320 3610
rect 6620 3430 9330 3640
rect 10330 3480 20840 3640
rect 10290 3460 20840 3480
rect 10120 3440 20840 3460
rect 10120 3420 10490 3440
rect 10290 3410 10420 3420
rect 12030 750 12220 3440
rect 13630 3430 20840 3440
<< viali >>
rect 830 5890 870 6050
rect 1010 5890 1050 6050
rect 730 5770 1050 5840
rect 830 5600 870 5710
rect 1110 5700 1190 5910
rect 810 4050 870 4230
rect 990 4050 1050 4230
rect 720 3940 1040 4000
rect 820 3760 860 3890
rect 1100 3870 1180 4070
<< metal1 >>
rect 1780 19890 18780 19950
rect 15580 19280 15710 19890
rect 15670 19050 15710 19280
rect 17330 19270 17480 19890
rect 17410 19050 17480 19270
rect 1430 18800 1440 18960
rect 1590 18800 1600 18960
rect 1440 14770 1590 18800
rect 15580 18780 15710 19050
rect 17330 18780 17480 19050
rect 1780 18720 18780 18780
rect 15580 16140 15710 18720
rect 15580 15760 15740 16140
rect 17330 15760 17480 18720
rect 1770 15700 18770 15760
rect 15580 15510 15740 15700
rect 15580 15090 15710 15510
rect 17330 15090 17480 15700
rect 15670 14860 15710 15090
rect 1430 14610 1440 14770
rect 1590 14610 1600 14770
rect 1440 10580 1590 14610
rect 15580 14590 15710 14860
rect 17410 14850 17480 15090
rect 17330 14590 17480 14850
rect 1770 14530 18770 14590
rect 1770 11730 1820 11840
rect 1430 10420 1440 10580
rect 1590 10420 1600 10580
rect 1770 10400 1820 11630
rect 15580 11570 15710 14530
rect 17330 11840 17480 14530
rect 17330 11740 17460 11840
rect 2600 11510 17270 11570
rect 17640 11510 18770 11570
rect 15580 10920 15710 11510
rect 15670 10670 15710 10920
rect 15580 10400 15710 10670
rect 1770 10340 17270 10400
rect 17720 10340 18770 10400
rect 1770 10130 1820 10340
rect 15580 7400 15710 10340
rect 17940 7520 17950 7620
rect 18210 7520 18220 7620
rect 19120 7610 19220 10650
rect 20800 10480 20810 10640
rect 20910 10480 20920 10640
rect 20510 10050 20640 10370
rect 20520 9760 20640 10050
rect 20810 9790 20910 10480
rect 20510 9190 20640 9760
rect 20520 8940 20640 9190
rect 20510 8780 20640 8940
rect 20520 8540 20640 8780
rect 20510 7920 20640 8540
rect 20520 7670 20640 7920
rect 19900 7580 20160 7660
rect 20510 7590 20640 7670
rect 20700 9640 20910 9790
rect 19900 7510 19920 7580
rect 20140 7510 20160 7580
rect 19900 7400 20160 7510
rect 15580 7310 20160 7400
rect 20700 7140 20810 9640
rect 2940 7090 6310 7120
rect 2940 6970 3400 7090
rect 3630 6970 4540 7090
rect 4770 6970 5540 7090
rect 5770 6970 6310 7090
rect 2940 6960 6310 6970
rect 6400 6990 9770 7100
rect 6400 6920 6710 6990
rect 3090 6750 6710 6920
rect 2840 6700 6100 6710
rect 2840 6510 2850 6700
rect 3020 6510 6100 6700
rect 2840 6500 6100 6510
rect 6400 6530 6710 6750
rect 2970 6420 6310 6440
rect 2970 6300 3130 6420
rect 3320 6300 3830 6420
rect 4020 6300 4980 6420
rect 5170 6300 6310 6420
rect 2970 6290 6310 6300
rect 6400 6360 9770 6530
rect 660 6230 6300 6240
rect 660 6120 1450 6230
rect 1680 6120 2350 6230
rect 2580 6120 3400 6230
rect 3630 6120 4540 6230
rect 660 6110 4540 6120
rect 4770 6110 5540 6230
rect 5770 6110 6300 6230
rect 660 6100 6300 6110
rect 824 6050 876 6062
rect 824 5890 830 6050
rect 870 5940 876 6050
rect 1004 6050 1056 6062
rect 2840 6050 2850 6070
rect 1004 5940 1010 6050
rect 870 5890 1010 5940
rect 1050 5940 1056 6050
rect 1050 5922 1190 5940
rect 1050 5910 1196 5922
rect 1050 5890 1110 5910
rect 824 5880 1110 5890
rect 824 5878 876 5880
rect 1004 5878 1056 5880
rect 718 5840 1062 5846
rect 718 5770 730 5840
rect 1050 5770 1062 5840
rect 718 5764 1062 5770
rect 824 5720 876 5722
rect 1104 5720 1110 5880
rect 824 5710 1110 5720
rect 824 5600 830 5710
rect 870 5700 1110 5710
rect 1190 5840 1196 5910
rect 1390 5890 2850 6050
rect 3020 5890 3030 6070
rect 6400 6050 6710 6360
rect 1390 5880 3030 5890
rect 3080 5890 6710 6050
rect 3080 5880 9770 5890
rect 1190 5780 2680 5840
rect 2840 5830 3030 5880
rect 1190 5700 1196 5780
rect 870 5688 1196 5700
rect 870 5660 1190 5688
rect 870 5600 876 5660
rect 2840 5640 6090 5830
rect 6400 5720 9770 5880
rect 824 5588 876 5600
rect 660 5540 6310 5560
rect 660 5400 700 5540
rect 920 5400 1820 5540
rect 2040 5400 3130 5540
rect 3320 5400 3830 5540
rect 4020 5520 6310 5540
rect 4020 5400 4980 5520
rect 5170 5400 6310 5520
rect 660 5390 6310 5400
rect 2960 5290 6290 5310
rect 2960 5160 3400 5290
rect 3630 5160 4540 5290
rect 2960 5150 4540 5160
rect 4770 5270 6290 5290
rect 4770 5150 5540 5270
rect 5770 5150 6290 5270
rect 2960 5140 6290 5150
rect 6400 5260 6710 5720
rect 6400 5150 9770 5260
rect 3080 5070 6170 5080
rect 3080 4920 5880 5070
rect 6160 4920 6170 5070
rect 6400 4960 6710 5150
rect 4260 4860 5820 4870
rect 2930 4850 5820 4860
rect 2850 4740 2860 4850
rect 2980 4740 5820 4850
rect 2930 4730 5820 4740
rect 6400 4850 9260 4960
rect 10180 4880 10490 7100
rect 15360 7030 20810 7140
rect 13800 6190 14180 6620
rect 14510 6190 14890 6620
rect 15360 6190 15490 7030
rect 15690 6180 16220 6650
rect 16060 5240 16220 6180
rect 16410 6170 16820 6630
rect 16060 5170 20880 5240
rect 20790 5010 20880 5170
rect 17390 4960 17540 5010
rect 20740 4960 20880 5010
rect 2960 4580 6290 4590
rect 2960 4570 3830 4580
rect 2960 4480 3130 4570
rect 3320 4480 3830 4570
rect 4020 4480 4980 4580
rect 5170 4480 6290 4580
rect 2960 4470 6290 4480
rect 650 4400 4540 4410
rect 650 4290 1450 4400
rect 1680 4390 3400 4400
rect 1680 4290 2350 4390
rect 2580 4290 3400 4390
rect 3630 4290 4540 4400
rect 4770 4290 5540 4410
rect 5770 4290 6320 4410
rect 650 4280 6320 4290
rect 6400 4390 6710 4850
rect 10170 4650 10180 4880
rect 10470 4650 10490 4880
rect 14460 4740 14470 4890
rect 14940 4840 14950 4890
rect 17390 4840 17480 4960
rect 14940 4740 17480 4840
rect 804 4230 876 4242
rect 804 4050 810 4230
rect 870 4110 876 4230
rect 984 4230 1056 4242
rect 984 4110 990 4230
rect 870 4050 990 4110
rect 1050 4110 1056 4230
rect 6400 4230 9170 4390
rect 3070 4200 6160 4210
rect 1370 4190 2980 4200
rect 1050 4082 1180 4110
rect 1050 4070 1186 4082
rect 1050 4050 1100 4070
rect 804 4040 1100 4050
rect 804 4038 876 4040
rect 984 4038 1056 4040
rect 510 4006 1050 4010
rect 510 4000 1052 4006
rect 510 3940 720 4000
rect 1040 3940 1052 4000
rect 510 3934 1052 3940
rect 510 3930 1050 3934
rect 814 3890 866 3902
rect 1094 3890 1100 4040
rect 1180 4000 1186 4070
rect 1370 4070 2870 4190
rect 2970 4070 2980 4190
rect 1370 4060 2980 4070
rect 1180 3980 2660 4000
rect 814 3760 820 3890
rect 860 3870 1100 3890
rect 860 3850 1110 3870
rect 1260 3850 2660 3980
rect 2860 3990 2980 4060
rect 3070 4050 5880 4200
rect 6160 4050 6170 4200
rect 2860 3850 6060 3990
rect 860 3840 2660 3850
rect 860 3760 866 3840
rect 1110 3830 2660 3840
rect 814 3748 866 3760
rect 6400 3770 6710 4230
rect 650 3580 700 3700
rect 920 3580 1820 3700
rect 2040 3580 3130 3700
rect 3320 3580 3830 3700
rect 4020 3580 4980 3700
rect 5170 3580 6320 3700
rect 6400 3660 9260 3770
rect 10180 3660 10490 4650
rect 14470 4190 14580 4740
rect 17390 4500 17480 4740
rect 20790 4500 20880 4960
rect 17390 4450 17550 4500
rect 20730 4450 20880 4500
rect 17390 4390 17480 4450
rect 20790 4390 20880 4450
rect 17390 4340 17550 4390
rect 20730 4340 20880 4390
rect 650 3570 6320 3580
rect 9850 3500 9860 3630
rect 10050 3590 10060 3630
rect 13790 3590 13880 4190
rect 14110 3750 14580 4190
rect 14810 3750 14820 3900
rect 14930 3750 14940 3900
rect 15390 3750 15820 4200
rect 16110 3750 16520 4210
rect 10050 3500 13880 3590
rect 16750 3660 16880 4200
rect 17390 3880 17480 4340
rect 20790 3880 20880 4340
rect 17390 3830 17550 3880
rect 20740 3830 20880 3880
rect 16750 3560 20840 3660
rect 200 3390 210 3470
rect 400 3390 410 3470
rect 20 3330 1450 3390
rect 20740 880 20840 3560
rect 20740 810 20960 880
rect 20 640 20150 690
rect 20 130 20150 180
rect 1760 -1670 1830 130
rect 1760 -1840 1810 -1670
rect 1760 -2780 1830 -1840
rect 3500 -2780 3570 130
rect 5240 -2780 5310 130
rect 6980 -2780 7050 130
rect 8720 -2780 8790 130
rect 10460 -2780 10530 130
rect 12200 -2780 12270 130
rect 13940 -2780 14010 130
rect 15680 -2780 15750 130
rect 17420 -2780 17490 130
rect 20890 70 20960 810
rect 20800 0 20810 70
rect 20960 0 20970 70
rect 1760 -2830 19010 -2780
rect 1760 -3290 1830 -2830
rect 3500 -3290 3570 -2830
rect 5240 -3290 5310 -2830
rect 6980 -3290 7050 -2830
rect 8720 -3290 8790 -2830
rect 10460 -3290 10530 -2830
rect 12200 -3290 12270 -2830
rect 13940 -3290 14010 -2830
rect 15680 -3290 15750 -2830
rect 17420 -3290 17490 -2830
rect 1760 -3340 19010 -3290
rect 1760 -5130 1830 -3340
rect 1760 -5340 1810 -5130
rect 1760 -5720 1830 -5340
rect 1760 -6030 1820 -5720
rect 1760 -6250 1830 -6030
rect 3500 -6250 3570 -3340
rect 5240 -6250 5310 -3340
rect 6980 -6250 7050 -3340
rect 8720 -6250 8790 -3340
rect 10460 -6250 10530 -3340
rect 12200 -6250 12270 -3340
rect 13940 -6250 14010 -3340
rect 15680 -6250 15750 -3340
rect 17420 -6250 17490 -3340
rect 1760 -6300 18850 -6250
rect 1760 -6760 1830 -6300
rect 3500 -6760 3570 -6300
rect 5240 -6760 5310 -6300
rect 6980 -6760 7050 -6300
rect 8720 -6760 8790 -6300
rect 10460 -6760 10530 -6300
rect 12200 -6760 12270 -6300
rect 13940 -6760 14010 -6300
rect 15680 -6760 15750 -6300
rect 17420 -6760 17490 -6300
rect 1760 -6810 18850 -6760
<< via1 >>
rect 1440 18800 1590 18960
rect 1440 14610 1590 14770
rect 1440 10420 1590 10580
rect 17950 7520 18210 7620
rect 20810 10480 20910 10640
rect 19920 7510 20140 7580
rect 3400 6970 3630 7090
rect 4540 6970 4770 7090
rect 5540 6970 5770 7090
rect 2850 6510 3020 6700
rect 3130 6300 3320 6420
rect 3830 6300 4020 6420
rect 4980 6300 5170 6420
rect 1450 6120 1680 6230
rect 2350 6120 2580 6230
rect 3400 6120 3630 6230
rect 4540 6110 4770 6230
rect 5540 6110 5770 6230
rect 730 5770 1050 5840
rect 2850 5890 3020 6070
rect 700 5400 920 5540
rect 1820 5400 2040 5540
rect 3130 5400 3320 5540
rect 3830 5400 4020 5540
rect 4980 5400 5170 5520
rect 3400 5160 3630 5290
rect 4540 5150 4770 5290
rect 5540 5150 5770 5270
rect 5880 4920 6160 5070
rect 2860 4740 2980 4850
rect 3130 4480 3320 4570
rect 3830 4480 4020 4580
rect 4980 4480 5170 4580
rect 1450 4290 1680 4400
rect 2350 4290 2580 4390
rect 3400 4290 3630 4400
rect 4540 4290 4770 4410
rect 5540 4290 5770 4410
rect 10180 4650 10470 4880
rect 14470 4740 14940 4890
rect 2870 4070 2970 4190
rect 1110 3870 1180 3980
rect 1180 3870 1260 3980
rect 1110 3850 1260 3870
rect 5880 4050 6160 4200
rect 700 3580 920 3700
rect 1820 3580 2040 3700
rect 3130 3580 3320 3700
rect 3830 3580 4020 3700
rect 4980 3580 5170 3700
rect 9860 3500 10050 3630
rect 14820 3750 14930 3900
rect 210 3390 400 3470
rect 20810 0 20960 70
<< metal2 >>
rect 1280 20070 1720 20080
rect 1720 20050 20470 20070
rect 1720 19710 19240 20050
rect 1720 19090 19240 19380
rect 20460 19710 20470 20050
rect 20460 19090 20470 19380
rect 1720 19080 20470 19090
rect 1280 19070 1720 19080
rect 1440 18960 1590 18970
rect 1590 18800 19010 18960
rect 1440 18790 1590 18800
rect 1730 17620 19030 18140
rect 1730 16610 19030 16870
rect 1730 15950 19030 16230
rect 1280 15880 1720 15890
rect 1720 15860 20470 15880
rect 1720 15520 19240 15860
rect 1720 15180 1780 15520
rect 1720 14900 19240 15180
rect 20460 15520 20470 15860
rect 20460 14900 20470 15180
rect 1720 14890 20470 14900
rect 1280 14880 1720 14890
rect 1440 14770 1590 14780
rect 1590 14610 19010 14770
rect 1440 14600 1590 14610
rect 1790 13430 19040 13950
rect 1730 12420 19030 12680
rect 19220 12240 20470 12270
rect 1730 11760 19030 12040
rect 19220 11740 19240 12240
rect 20460 11740 20470 12240
rect 1290 11660 1720 11670
rect 1280 11330 1290 11610
rect 1280 10710 1290 10970
rect 19220 11610 20470 11740
rect 1720 11330 20770 11610
rect 1720 10710 20770 10970
rect 1280 10700 20770 10710
rect 20810 10640 20910 10850
rect 1440 10580 1590 10590
rect 1590 10420 17240 10580
rect 17720 10440 19000 10580
rect 20810 10470 20910 10480
rect 17720 10420 18880 10440
rect 1440 10410 1590 10420
rect 1800 9240 17290 9760
rect 1800 8230 17290 8490
rect 1800 7490 17290 7850
rect 17950 7620 18210 7630
rect 17950 7510 18210 7520
rect 19900 7580 20160 7760
rect 19900 7510 19920 7580
rect 20140 7510 20160 7580
rect 19900 7490 20160 7510
rect 8300 7260 12010 7270
rect 1450 7250 1680 7260
rect 1450 6230 1680 7000
rect 730 5840 1050 5850
rect 1050 5770 1260 5840
rect 730 5710 1260 5770
rect 700 5540 920 5560
rect 700 3710 920 5400
rect 1110 3980 1260 5710
rect 1450 4400 1680 6120
rect 2350 7250 2580 7260
rect 2350 6230 2580 7000
rect 3400 7250 3630 7260
rect 1450 4280 1680 4290
rect 1820 5540 2040 5560
rect 1110 3840 1260 3850
rect 70 3470 560 3610
rect 700 3560 920 3570
rect 1820 3700 2040 5400
rect 2350 4390 2580 6120
rect 2840 6700 3030 6710
rect 2840 6510 2850 6700
rect 3020 6510 3030 6700
rect 2840 6070 3030 6510
rect 2840 5890 2850 6070
rect 3020 5890 3030 6070
rect 2840 5880 3030 5890
rect 3130 6420 3320 6440
rect 3130 5540 3320 6300
rect 2350 4280 2580 4290
rect 2860 4850 2980 4860
rect 2860 4190 2980 4740
rect 2860 4070 2870 4190
rect 2970 4070 2980 4190
rect 3130 4570 3320 5400
rect 2870 4060 2970 4070
rect 1820 3550 2040 3560
rect 3130 3700 3320 4480
rect 3400 6230 3630 6970
rect 4540 7250 4770 7260
rect 3400 5290 3630 6120
rect 3400 4400 3630 5160
rect 3400 4280 3630 4290
rect 3830 6420 4020 6440
rect 3830 5540 4020 6300
rect 3830 4580 4020 5400
rect 3130 3550 3320 3560
rect 3830 3700 4020 4480
rect 4540 6230 4770 6970
rect 5540 7250 5770 7260
rect 4540 5290 4770 6110
rect 4540 4410 4770 5150
rect 4540 4280 4770 4290
rect 4980 6420 5170 6440
rect 4980 5520 5170 6300
rect 4980 4580 5170 5400
rect 3830 3550 4020 3560
rect 4980 3700 5170 4480
rect 5540 6230 5770 6970
rect 6850 6830 8300 7210
rect 12010 6830 13380 7210
rect 6850 6810 13380 6830
rect 6750 6680 9700 6710
rect 6750 6220 6800 6680
rect 8210 6220 9700 6680
rect 6750 6180 9700 6220
rect 10530 6180 14460 6710
rect 5540 5270 5770 6110
rect 6850 6060 13380 6080
rect 6850 5560 8300 6060
rect 12010 5560 13380 6060
rect 6850 5540 13380 5560
rect 13570 5440 14460 6180
rect 5540 4410 5770 5150
rect 6760 5420 10050 5440
rect 5540 4280 5770 4290
rect 5870 5070 6170 5080
rect 5870 4920 5880 5070
rect 6160 4920 6170 5070
rect 5870 4870 6170 4920
rect 5870 4660 5880 4870
rect 6160 4660 6170 4870
rect 6760 4970 6800 5420
rect 10010 4970 10050 5420
rect 6760 4670 10050 4970
rect 10530 5090 14460 5440
rect 18640 5110 19600 5120
rect 5870 4200 6170 4660
rect 5870 4050 5880 4200
rect 6160 4050 6170 4200
rect 6760 4550 9170 4560
rect 5880 4040 6160 4050
rect 6760 4040 9170 4050
rect 9280 3950 10050 4670
rect 10180 4880 10470 4890
rect 10530 4670 13210 5090
rect 10180 4640 10470 4650
rect 10530 4550 13000 4560
rect 10530 4040 13000 4050
rect 13060 3950 13210 4670
rect 4980 3550 5170 3560
rect 6750 3630 10050 3950
rect 6750 3550 9860 3630
rect 10540 3760 13210 3950
rect 14220 5060 14460 5090
rect 14220 3760 14360 5060
rect 14470 4890 14940 4900
rect 17640 4800 18640 5110
rect 19600 4930 20620 5110
rect 19600 4800 20630 4930
rect 17640 4780 20630 4800
rect 14470 4730 14940 4740
rect 17530 4640 19020 4670
rect 18500 4200 19020 4640
rect 17530 4160 19020 4200
rect 19260 4630 20750 4670
rect 19260 4190 19700 4630
rect 20670 4190 20750 4630
rect 19260 4160 20750 4190
rect 17470 4040 20750 4050
rect 10540 3660 14360 3760
rect 14820 3900 14930 3910
rect 14820 3740 14930 3750
rect 14830 3660 14920 3740
rect 10540 3550 14920 3660
rect 17470 3730 18640 4040
rect 19600 3730 20750 4040
rect 9860 3490 10050 3500
rect 70 3390 210 3470
rect 400 3390 560 3470
rect 70 3320 560 3390
rect 1810 3120 16900 3460
rect 17470 3120 20750 3730
rect 1810 2510 16900 2730
rect 17470 2510 20380 2730
rect 1810 1890 16900 2110
rect 17470 1890 20380 2110
rect 1810 1270 16900 1490
rect 17470 1270 20380 1490
rect 3550 1170 3620 1200
rect 5290 1170 5360 1200
rect 6950 1170 7100 1200
rect 8760 1170 8890 1200
rect 10500 1170 10630 1200
rect 12240 1170 12320 1200
rect 13970 1170 14070 1200
rect 15720 1170 15820 1200
rect 1870 1140 17000 1170
rect 1870 1020 1890 1140
rect 2040 1020 17000 1140
rect 1890 990 2040 1000
rect 18900 460 19340 600
rect 130 350 20750 360
rect 20750 340 20790 350
rect 20790 70 20960 80
rect 20790 0 20810 70
rect 20790 -10 20960 0
rect 130 -40 19240 -30
rect 19240 -50 20790 -40
rect 1810 -350 18640 -120
rect 1810 -960 18640 -740
rect 1810 -1580 18640 -1360
rect 2170 -1830 18750 -1680
rect 1810 -2200 18640 -1980
rect 1880 -2310 2090 -2300
rect 1880 -2520 2090 -2510
rect 130 -2910 1680 -2900
rect 19240 -2940 20790 -2930
rect 1680 -3110 19240 -3100
rect 1680 -3500 19240 -3490
rect 1810 -3820 18640 -3600
rect 130 -3960 1680 -3950
rect 19240 -3990 20790 -3980
rect 1810 -4430 18640 -4210
rect 1810 -5050 18640 -4830
rect 2920 -5300 18750 -5150
rect 1810 -5670 18640 -5450
rect 1880 -5790 2040 -5780
rect 130 -5930 1680 -5920
rect 120 -6590 130 -6580
rect 1880 -5970 2040 -5960
rect 19240 -5940 20790 -5930
rect 1680 -6590 19240 -6580
rect 120 -6980 19240 -6970
rect 19240 -6990 20790 -6980
<< via2 >>
rect 1280 19080 1720 20070
rect 19240 19090 20460 20050
rect 1280 14890 1720 15880
rect 19240 14900 20460 15860
rect 19240 11740 20460 12240
rect 1290 10710 1720 11660
rect 17950 7520 18210 7620
rect 1450 7000 1680 7250
rect 2350 7000 2580 7250
rect 3400 7090 3630 7250
rect 3400 7000 3630 7090
rect 700 3700 920 3710
rect 700 3580 920 3700
rect 700 3570 920 3580
rect 1820 3580 2040 3700
rect 1820 3560 2040 3580
rect 4540 7090 4770 7250
rect 4540 7000 4770 7090
rect 3130 3580 3320 3700
rect 3130 3560 3320 3580
rect 5540 7090 5770 7250
rect 5540 7000 5770 7090
rect 3830 3580 4020 3700
rect 3830 3560 4020 3580
rect 8300 6830 12010 7260
rect 6800 6220 8210 6680
rect 8300 5560 12010 6060
rect 5880 4660 6160 4870
rect 6800 4970 10010 5420
rect 6760 4050 9170 4550
rect 10180 4650 10470 4880
rect 10530 4050 13000 4550
rect 4980 3580 5170 3700
rect 4980 3560 5170 3580
rect 13210 3760 14220 5090
rect 14470 4740 14940 4890
rect 18640 4800 19600 5110
rect 17530 4200 18500 4640
rect 19700 4190 20670 4630
rect 18640 3730 19600 4040
rect 1890 1000 2040 1140
rect 130 340 20750 350
rect 130 -30 20790 340
rect 19240 -40 20790 -30
rect 1880 -2510 2090 -2310
rect 130 -3110 1680 -2910
rect 19240 -3110 20790 -2940
rect 130 -3490 20790 -3110
rect 130 -3950 1680 -3490
rect 19240 -3980 20790 -3490
rect 130 -6590 1680 -5930
rect 1880 -5960 2040 -5790
rect 19240 -6590 20790 -5940
rect 120 -6970 20790 -6590
rect 19240 -6980 20790 -6970
<< metal3 >>
rect 1270 20070 1730 20075
rect 1270 19080 1280 20070
rect 2200 20040 2210 20070
rect 19230 20050 20470 20055
rect 19230 20040 19240 20050
rect 2200 19720 19240 20040
rect 2200 19080 2210 19720
rect 19230 19090 19240 19720
rect 20460 19090 20470 20050
rect 19230 19085 20470 19090
rect 1270 19075 1730 19080
rect 9390 18600 12140 18960
rect 9900 17630 9910 18130
rect 10920 17630 10930 18130
rect 9900 16610 9910 16870
rect 10920 16610 10930 16870
rect 9390 15960 9400 16230
rect 11920 15960 11930 16230
rect 1270 15880 1730 15885
rect 1270 14880 1280 15880
rect 1720 15870 1730 15880
rect 2200 15850 2210 15870
rect 19230 15860 20470 15865
rect 19230 15850 19240 15860
rect 2200 15530 19240 15850
rect 2200 14880 2210 15530
rect 19230 14900 19240 15530
rect 20460 14900 20470 15860
rect 19230 14895 20470 14900
rect 9390 14410 12140 14770
rect 9900 13440 9910 13940
rect 10920 13440 10930 13940
rect 9900 12420 9910 12680
rect 10920 12420 10930 12680
rect 19230 12240 20470 12245
rect 9390 11760 9400 12030
rect 11920 11760 11930 12030
rect 19230 11740 19240 12240
rect 20460 11740 20470 12240
rect 19230 11735 20470 11740
rect 1710 11665 1810 11670
rect 1280 11660 1810 11665
rect 1280 10710 1290 11660
rect 1720 11650 19230 11660
rect 2200 11340 19230 11650
rect 2200 10790 2210 11340
rect 2200 10710 2230 10790
rect 1280 10705 2230 10710
rect 1700 10700 2230 10705
rect 9390 10220 12140 10580
rect 19220 10370 19230 11340
rect 19600 11340 20360 11660
rect 19600 10370 19610 11340
rect 20350 10370 20360 11340
rect 20760 10370 20770 11660
rect 9900 9250 9910 9750
rect 10920 9250 10930 9750
rect 9900 8230 9910 8490
rect 10920 8230 10930 8490
rect 9390 7490 9400 7850
rect 12130 7490 12140 7850
rect 17460 7650 19030 7840
rect 17430 7620 19050 7650
rect 17430 7520 17950 7620
rect 18210 7520 19050 7620
rect 1340 6990 1350 7290
rect 1940 7255 5770 7290
rect 8290 7260 12020 7265
rect 1940 7250 5780 7255
rect 1940 7000 2350 7250
rect 2580 7000 3400 7250
rect 3630 7000 4540 7250
rect 4770 7000 5540 7250
rect 5770 7000 5780 7250
rect 1940 6995 5780 7000
rect 1940 6990 5770 6995
rect 8290 6830 8300 7260
rect 12010 6830 12020 7260
rect 17430 7240 19050 7520
rect 8290 6825 9430 6830
rect 6790 6680 8220 6685
rect 6790 6220 6800 6680
rect 8210 6220 8220 6680
rect 6790 6215 8220 6220
rect 6800 5425 8210 6215
rect 8300 6065 9430 6825
rect 8290 6060 9430 6065
rect 11980 6825 12020 6830
rect 11980 6065 12010 6825
rect 11980 6060 12020 6065
rect 8290 5560 8300 6060
rect 12010 5560 12020 6060
rect 8290 5555 12020 5560
rect 8300 5540 12010 5555
rect 6790 5420 10020 5425
rect 6780 4970 6790 5420
rect 10010 4970 10020 5420
rect 6790 4965 10020 4970
rect 13200 5090 14230 5095
rect 5830 4880 6170 4885
rect 10170 4880 10480 4885
rect 5830 4870 10180 4880
rect 5830 4660 5880 4870
rect 6160 4660 10180 4870
rect 5830 4650 10180 4660
rect 10470 4840 10480 4880
rect 10470 4650 10490 4840
rect 5830 4645 6170 4650
rect 10170 4645 10480 4650
rect 7710 4555 11940 4560
rect 6750 4550 13010 4555
rect 6750 4050 6760 4550
rect 9170 4050 9340 4550
rect 13000 4050 13010 4550
rect 6750 4045 13010 4050
rect 7710 4040 11940 4045
rect 680 3560 690 3830
rect 1250 3705 5170 3830
rect 13200 3760 13210 5090
rect 14220 3760 14230 5090
rect 14460 4890 14950 4895
rect 14460 4740 14470 4890
rect 14940 4740 14950 4890
rect 14460 4735 14950 4740
rect 17540 4645 18510 7240
rect 19200 7230 20770 7840
rect 18630 5110 19610 5115
rect 18630 4800 18640 5110
rect 19600 4800 19610 5110
rect 18630 4795 19610 4800
rect 17520 4640 18510 4645
rect 17520 4200 17530 4640
rect 18500 4200 18510 4640
rect 17520 4195 18510 4200
rect 17540 4190 18510 4195
rect 18640 4045 19600 4795
rect 19700 4635 20670 7230
rect 19690 4630 20680 4635
rect 19690 4190 19700 4630
rect 20670 4190 20680 4630
rect 19690 4185 20680 4190
rect 13200 3755 14230 3760
rect 18630 4040 19610 4045
rect 18630 3730 18640 4040
rect 19600 3730 19610 4040
rect 18630 3725 19610 3730
rect 1250 3700 5180 3705
rect 1250 3560 1820 3700
rect 2040 3560 3130 3700
rect 3320 3560 3830 3700
rect 4020 3560 4980 3700
rect 5170 3560 5180 3700
rect 1810 3555 2050 3560
rect 3120 3555 3330 3560
rect 3820 3555 4030 3560
rect 4970 3555 5180 3560
rect 1800 3300 16900 3460
rect 1800 3120 8770 3300
rect 8760 1270 8770 3120
rect 9460 3120 10510 3300
rect 9460 1270 9470 3120
rect 10500 1270 10510 3120
rect 11200 3120 16900 3300
rect 11200 1270 11210 3120
rect 1880 1140 2050 1145
rect 1880 1000 1890 1140
rect 2040 1000 2050 1140
rect 1880 995 2050 1000
rect 19240 590 20780 600
rect 130 360 20780 590
rect 120 350 20780 360
rect 120 -700 130 350
rect 20750 345 20780 350
rect 20750 340 20800 345
rect 1680 -35 19240 -30
rect 1680 -700 1690 -35
rect 1810 -170 18640 -120
rect 1810 -350 8770 -170
rect 120 -705 1690 -700
rect 8760 -2200 8770 -350
rect 9460 -350 10510 -170
rect 9460 -2200 9470 -350
rect 10500 -2200 10510 -350
rect 11200 -350 18640 -170
rect 11200 -2200 11210 -350
rect 19230 -700 19240 -35
rect 20790 -700 20800 340
rect 19230 -705 20800 -700
rect 1870 -2310 2100 -2305
rect 1870 -2510 1880 -2310
rect 2090 -2510 2100 -2310
rect 1870 -2515 2100 -2510
rect 130 -2905 20790 -2860
rect 120 -2910 20790 -2905
rect 120 -3950 130 -2910
rect 1680 -2935 20790 -2910
rect 1680 -2940 20800 -2935
rect 1680 -3110 19240 -2940
rect 1680 -3495 19240 -3490
rect 1680 -3950 1690 -3495
rect 1810 -3820 8770 -3600
rect 120 -3955 1690 -3950
rect 8760 -5670 8770 -3820
rect 9460 -3820 10490 -3600
rect 9460 -5670 9470 -3820
rect 10480 -5670 10490 -3820
rect 11190 -3820 18640 -3600
rect 11190 -5670 11200 -3820
rect 19230 -3980 19240 -3495
rect 20790 -3980 20800 -2940
rect 19230 -3985 20800 -3980
rect 1870 -5790 2050 -5785
rect 120 -5930 1690 -5925
rect 120 -6585 130 -5930
rect 110 -6590 130 -6585
rect 110 -6970 120 -6590
rect 1680 -6350 1690 -5930
rect 1870 -5960 1880 -5790
rect 2040 -5960 2050 -5790
rect 1870 -5965 2050 -5960
rect 19230 -5940 20800 -5935
rect 19230 -6350 19240 -5940
rect 1680 -6590 19240 -6350
rect 110 -6975 19240 -6970
rect 19230 -6980 19240 -6975
rect 20790 -6980 20800 -5940
rect 19230 -6985 20800 -6980
<< via3 >>
rect 1280 19080 1720 20070
rect 1720 19080 2200 20070
rect 19240 19090 20460 20050
rect 9910 17630 10920 18130
rect 9910 16610 10920 16870
rect 9400 15960 11920 16230
rect 1280 14890 1720 15870
rect 1720 14890 2200 15870
rect 1280 14880 2200 14890
rect 19240 14900 20460 15860
rect 9910 13440 10920 13940
rect 9910 12420 10920 12680
rect 9400 11760 11920 12030
rect 19240 11740 20460 12240
rect 1290 10710 1720 11650
rect 1720 10710 2200 11650
rect 19230 10370 19600 11660
rect 20360 10370 20760 11660
rect 9910 9250 10920 9750
rect 9910 8230 10920 8490
rect 9400 7490 12130 7850
rect 1350 7250 1940 7290
rect 1350 7000 1450 7250
rect 1450 7000 1680 7250
rect 1680 7000 1940 7250
rect 1350 6990 1940 7000
rect 9430 6830 11980 7230
rect 9430 6060 11980 6830
rect 9430 5610 11980 6060
rect 6790 4970 6800 5420
rect 6800 4970 10010 5420
rect 9340 4050 10530 4550
rect 10530 4050 12130 4550
rect 690 3710 1250 3830
rect 690 3570 700 3710
rect 700 3570 920 3710
rect 920 3570 1250 3710
rect 13210 3760 14220 5090
rect 14470 4740 14940 4890
rect 690 3560 1250 3570
rect 8770 1270 9460 3300
rect 10510 1270 11200 3300
rect 1890 1000 2040 1130
rect 130 -30 1680 350
rect 130 -700 1680 -30
rect 8770 -2200 9460 -170
rect 10510 -2200 11200 -170
rect 19240 -40 20790 340
rect 19240 -700 20790 -40
rect 1880 -2510 2090 -2310
rect 130 -3950 1680 -2910
rect 8770 -5670 9460 -3600
rect 10490 -5670 11190 -3600
rect 19240 -3980 20790 -2940
rect 130 -6970 1680 -5930
rect 1880 -5960 2040 -5790
rect 19240 -6980 20790 -5940
<< metal4 >>
rect 1279 19080 1280 20071
rect 2510 19090 2520 20090
rect 2200 19080 2520 19090
rect 1279 19079 2520 19080
rect 1280 15871 2520 19079
rect 19230 19090 19240 20090
rect 9400 18130 11910 18140
rect 9400 17630 9910 18130
rect 10920 17630 11910 18130
rect 9400 16870 11910 17630
rect 9400 16610 9910 16870
rect 10920 16610 11910 16870
rect 9400 16231 11910 16610
rect 9399 16230 11921 16231
rect 9399 15960 9400 16230
rect 11920 15960 12130 16230
rect 9399 15959 12130 15960
rect 1279 15870 2520 15871
rect 1279 14880 1280 15870
rect 2200 14880 2520 15870
rect 1279 14879 2520 14880
rect 1280 11650 2520 14879
rect 9400 14820 12130 15959
rect 19230 15860 20470 19090
rect 19230 14900 19240 15860
rect 20460 14900 20470 15860
rect 9400 14400 11920 14820
rect 9400 13940 12130 14400
rect 9400 13440 9910 13940
rect 10920 13440 12130 13940
rect 9400 12680 12130 13440
rect 9400 12420 9910 12680
rect 10920 12420 12130 12680
rect 9400 12031 12130 12420
rect 9399 12030 12130 12031
rect 9399 11760 9400 12030
rect 11920 11760 12130 12030
rect 9399 11759 12130 11760
rect 1280 10710 1290 11650
rect 2200 10710 2520 11650
rect 1280 7480 2520 10710
rect 9400 10680 12130 11759
rect 19230 12240 20470 14900
rect 19230 11740 19240 12240
rect 20460 11740 20470 12240
rect 19230 11661 20470 11740
rect 19229 11660 20761 11661
rect 9400 10080 11920 10680
rect 19229 10370 19230 11660
rect 19600 10370 20360 11660
rect 20760 10370 20761 11660
rect 19229 10369 20761 10370
rect 19230 10190 20470 10369
rect 9400 9750 12130 10080
rect 9400 9250 9910 9750
rect 10920 9250 12130 9750
rect 9400 8490 12130 9250
rect 9400 8230 9910 8490
rect 10920 8230 12130 8490
rect 9400 7851 12130 8230
rect 9399 7850 12131 7851
rect 9399 7490 9400 7850
rect 12130 7490 12131 7850
rect 9399 7489 12131 7490
rect 1350 7291 1940 7480
rect 1349 7290 1941 7291
rect 1349 6990 1350 7290
rect 1940 6990 1941 7290
rect 1349 6989 1941 6990
rect 9400 7230 12130 7489
rect 9400 5610 9430 7230
rect 11980 5610 12130 7230
rect 9400 5560 12130 5610
rect 6789 5420 10011 5421
rect 6789 4970 6790 5420
rect 10010 4970 10011 5420
rect 6789 4969 10011 4970
rect 13209 5090 14221 5091
rect 9340 4551 12140 4570
rect 9339 4550 12140 4551
rect 9339 4050 9340 4550
rect 12130 4050 12140 4550
rect 9339 4049 12140 4050
rect 689 3830 1251 3831
rect 689 3560 690 3830
rect 1250 3560 1251 3830
rect 689 3559 1251 3560
rect 690 3440 1250 3559
rect 130 351 1680 3440
rect 9340 3301 12140 4049
rect 13209 3760 13210 5090
rect 14220 3760 14221 5090
rect 14470 4891 14940 5580
rect 14469 4890 14941 4891
rect 14469 4740 14470 4890
rect 14940 4740 14941 4890
rect 14469 4739 14941 4740
rect 13209 3759 14221 3760
rect 8769 3300 12140 3301
rect 8769 1270 8770 3300
rect 9460 1270 10510 3300
rect 11200 1270 12140 3300
rect 8769 1269 12140 1270
rect 1880 1130 2050 1140
rect 1880 1000 1890 1130
rect 2040 1000 2050 1130
rect 129 350 1681 351
rect 129 -700 130 350
rect 1680 -700 1681 350
rect 129 -701 1681 -700
rect 130 -2909 1680 -701
rect 1880 -2309 2050 1000
rect 9340 -169 12140 1269
rect 19240 341 20790 3430
rect 8769 -170 12140 -169
rect 8769 -2200 8770 -170
rect 9460 -2200 10510 -170
rect 11200 -2200 12140 -170
rect 19239 340 20791 341
rect 19239 -700 19240 340
rect 20790 -700 20791 340
rect 19239 -701 20791 -700
rect 8769 -2201 12140 -2200
rect 1879 -2310 2091 -2309
rect 1879 -2510 1880 -2310
rect 2090 -2510 2091 -2310
rect 1879 -2511 2091 -2510
rect 129 -2910 1681 -2909
rect 129 -3950 130 -2910
rect 1680 -3950 1681 -2910
rect 129 -3951 1681 -3950
rect 130 -5190 1680 -3951
rect 1650 -5929 1680 -5190
rect 1880 -5789 2050 -2511
rect 9340 -3599 12140 -2201
rect 19240 -2939 20790 -701
rect 8769 -3600 12140 -3599
rect 8769 -5670 8770 -3600
rect 9460 -5670 10490 -3600
rect 11190 -5670 12140 -3600
rect 19239 -2940 20791 -2939
rect 19239 -3980 19240 -2940
rect 20790 -3980 20791 -2940
rect 19239 -3981 20791 -3980
rect 8769 -5671 12140 -5670
rect 1879 -5790 2050 -5789
rect 1650 -5930 1681 -5929
rect 1680 -6970 1681 -5930
rect 1879 -5960 1880 -5790
rect 2040 -5960 2050 -5790
rect 1879 -5961 2041 -5960
rect 9340 -6040 12140 -5671
rect 19240 -5190 20790 -3981
rect 19240 -5939 19260 -5190
rect 19239 -5940 19260 -5939
rect 129 -6971 1681 -6970
rect 19239 -6980 19240 -5940
rect 20790 -6980 20791 -5939
rect 19239 -6981 20791 -6980
<< via4 >>
rect 1280 20070 2510 20090
rect 1280 19090 2200 20070
rect 2200 19090 2510 20070
rect 19240 20050 20470 20090
rect 19240 19090 20460 20050
rect 20460 19090 20470 20050
rect 6790 4970 10010 5420
rect 13210 3760 14220 4570
rect 120 -5930 1650 -5190
rect 120 -6970 130 -5930
rect 130 -6970 1650 -5930
rect 19260 -5940 20790 -5190
rect 19260 -6970 20790 -5940
<< metal5 >>
rect 1256 20100 2534 20114
rect 19216 20100 20494 20114
rect 1256 20090 20494 20100
rect 1256 19090 1280 20090
rect 2510 19430 19240 20090
rect 2510 19090 2534 19430
rect 1256 19066 2534 19090
rect 19216 19090 19240 19430
rect 20470 19090 20494 20090
rect 19216 19066 20494 19090
rect 1570 16080 2350 18340
rect 1570 15500 18420 16080
rect 1570 -5166 2350 15500
rect 6766 5440 10034 5444
rect 6766 5420 21080 5440
rect 6766 4970 6790 5420
rect 10010 4970 21080 5420
rect 6766 4946 21080 4970
rect 9850 4940 21080 4946
rect 13210 4594 21080 4610
rect 13186 4570 21080 4594
rect 13186 3760 13210 4570
rect 14220 4110 21080 4570
rect 14220 3760 14244 4110
rect 13186 3736 14244 3760
rect 96 -5190 2350 -5166
rect 96 -6970 120 -5190
rect 1650 -5830 2350 -5190
rect 19236 -5190 20814 -5166
rect 19236 -5830 19260 -5190
rect 1650 -6970 19260 -5830
rect 20790 -6970 20814 -5190
rect 96 -6980 20814 -6970
rect 96 -6994 1674 -6980
rect 19236 -6994 20814 -6980
use lvds_currm_n  lvds_currm_n_0
timestamp 1654683408
transform 1 0 140 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_1
timestamp 1654683408
transform 1 0 1880 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_2
timestamp 1654683408
transform 1 0 3620 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_3
timestamp 1654683408
transform 1 0 5360 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_4
timestamp 1654683408
transform 1 0 7100 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_5
timestamp 1654683408
transform 1 0 14060 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_6
timestamp 1654683408
transform 1 0 12320 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_7
timestamp 1654683408
transform 1 0 10580 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_8
timestamp 1654683408
transform 1 0 8840 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_9
timestamp 1654683408
transform 1 0 19280 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_10
timestamp 1654683408
transform 1 0 17540 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_11
timestamp 1654683408
transform 1 0 15800 0 1 600
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_12
timestamp 1654683408
transform 1 0 3620 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_13
timestamp 1654683408
transform 1 0 1880 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_14
timestamp 1654683408
transform 1 0 5360 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_15
timestamp 1654683408
transform 1 0 7100 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_16
timestamp 1654683408
transform 1 0 8840 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_17
timestamp 1654683408
transform 1 0 10580 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_18
timestamp 1654683408
transform 1 0 12320 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_19
timestamp 1654683408
transform 1 0 14060 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_20
timestamp 1654683408
transform 1 0 15800 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_21
timestamp 1654683408
transform 1 0 17540 0 1 -2870
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_22
timestamp 1654683408
transform 1 0 3620 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_23
timestamp 1654683408
transform 1 0 1880 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_24
timestamp 1654683408
transform 1 0 5360 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_25
timestamp 1654683408
transform 1 0 7100 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_26
timestamp 1654683408
transform 1 0 8840 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_27
timestamp 1654683408
transform 1 0 10580 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_28
timestamp 1654683408
transform 1 0 12320 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_29
timestamp 1654683408
transform 1 0 14060 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_30
timestamp 1654683408
transform 1 0 15800 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_n  lvds_currm_n_31
timestamp 1654683408
transform 1 0 17540 0 1 -6340
box -150 -600 1600 2884
use lvds_currm_p  lvds_currm_p_0
timestamp 1654683408
transform 1 0 3540 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_1
timestamp 1654683408
transform 1 0 1800 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_2
timestamp 1654683408
transform 1 0 5280 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_3
timestamp 1654683408
transform 1 0 7020 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_4
timestamp 1654683408
transform 1 0 8760 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_5
timestamp 1654683408
transform 1 0 17460 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_6
timestamp 1654683408
transform 1 0 15720 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_7
timestamp 1654683408
transform 1 0 13980 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_8
timestamp 1654683408
transform 1 0 12240 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_9
timestamp 1654683408
transform 1 0 10500 0 1 7500
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_10
timestamp 1654683408
transform 1 0 3540 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_11
timestamp 1654683408
transform 1 0 1800 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_12
timestamp 1654683408
transform 1 0 5280 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_13
timestamp 1654683408
transform 1 0 7020 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_14
timestamp 1654683408
transform 1 0 8760 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_15
timestamp 1654683408
transform 1 0 10500 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_16
timestamp 1654683408
transform 1 0 12240 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_17
timestamp 1654683408
transform 1 0 13980 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_18
timestamp 1654683408
transform 1 0 15720 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_19
timestamp 1654683408
transform 1 0 17460 0 1 11690
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_20
timestamp 1654683408
transform 1 0 3540 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_21
timestamp 1654683408
transform 1 0 1800 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_22
timestamp 1654683408
transform 1 0 5280 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_23
timestamp 1654683408
transform 1 0 7020 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_24
timestamp 1654683408
transform 1 0 8760 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_25
timestamp 1654683408
transform 1 0 10500 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_26
timestamp 1654683408
transform 1 0 12240 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_27
timestamp 1654683408
transform 1 0 13980 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_28
timestamp 1654683408
transform 1 0 15720 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_29
timestamp 1654683408
transform 1 0 17460 0 1 15880
box -70 -10 1680 4194
use lvds_currm_p  lvds_currm_p_30
timestamp 1654683408
transform 1 0 19200 0 1 7500
box -70 -10 1680 4194
use lvds_diffamp  lvds_diffamp_0
timestamp 1654683408
transform 1 0 17450 0 1 3750
box -60 -50 1690 1388
use lvds_diffamp  lvds_diffamp_1
timestamp 1654683408
transform 1 0 19190 0 1 3750
box -60 -50 1690 1388
use lvds_nswitch  lvds_nswitch_0
timestamp 1654683408
transform 1 0 6720 0 1 3690
box -100 -100 2634 1338
use lvds_nswitch  lvds_nswitch_1
timestamp 1654683408
transform 1 0 10500 0 1 3690
box -100 -100 2634 1338
use lvds_switch_p  lvds_switch_p_0
timestamp 1654683408
transform 1 0 6572 0 1 5076
box 48 -6 3262 2104
use lvds_switch_p  lvds_switch_p_1
timestamp 1654683408
transform 1 0 10352 0 1 5076
box 48 -6 3262 2104
use sky130_fd_pr__cap_mim_m3_1_N3PKNJ  sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0
timestamp 1654683408
transform -1 0 15679 0 -1 6300
box -3150 -1100 3149 1100
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#3  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1654683408
transform 0 -1 5991 1 0 16351
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#3  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_1
timestamp 1654683408
transform 0 -1 15641 1 0 16351
box -3351 -3101 3373 3101
use sky130_fd_pr__res_xhigh_po_0p35_RS2YEK  sky130_fd_pr__res_xhigh_po_0p35_RS2YEK_0
timestamp 1654683408
transform 1 0 16469 0 1 5188
box -519 -1598 519 1598
use sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL  sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL_0
timestamp 1654683408
transform 1 0 13990 0 1 5188
box -360 -1598 360 1598
use sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL  sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL_1
timestamp 1654683408
transform 1 0 14700 0 1 5188
box -360 -1598 360 1598
use sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL  sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL_2
timestamp 1654683408
transform 1 0 15600 0 1 5188
box -360 -1598 360 1598
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_0
timestamp 1649384327
transform 1 0 688 0 1 3659
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_1
timestamp 1649384327
transform 1 0 698 0 1 5489
box -38 -49 518 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_0
timestamp 1649384327
transform 1 0 1248 0 1 3659
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_1
timestamp 1649384327
transform 1 0 2948 0 1 3659
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_2
timestamp 1649384327
transform 1 0 4648 0 1 3659
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_3
timestamp 1649384327
transform 1 0 2958 0 1 4529
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_4
timestamp 1649384327
transform 1 0 4658 0 1 4529
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_5
timestamp 1649384327
transform 1 0 4678 0 1 6359
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_6
timestamp 1649384327
transform 1 0 4668 0 1 5489
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_7
timestamp 1649384327
transform 1 0 2978 0 1 6359
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_8
timestamp 1649384327
transform 1 0 1268 0 1 5489
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_9
timestamp 1649384327
transform 1 0 2968 0 1 5489
box -38 -49 1670 715
<< labels >>
rlabel metal5 1360 19290 1670 19720 1 VP
rlabel metal5 380 -6870 690 -6440 1 VN
rlabel metal1 510 3930 610 4010 1 In
rlabel metal5 20910 4160 21040 4580 1 OutP
rlabel metal5 20910 4960 21040 5380 1 OutN
rlabel metal4 10230 7330 10690 7430 1 vm6d
rlabel metal4 9890 3670 10350 3770 1 vm1d
rlabel metal1 6480 4080 6610 4230 1 vm2g
rlabel metal1 10210 4590 10340 4740 1 vm5g
rlabel metal1 17120 4750 17220 4830 1 vm20g
rlabel metal2 1130 4640 1230 4760 1 vx9y
rlabel metal1 1280 5780 1340 5810 1 vx14y
rlabel metal1 2890 5730 2990 5790 1 vx1y
rlabel metal1 2880 3870 2930 3960 1 vx6y
<< end >>
