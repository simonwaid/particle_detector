magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< pwell >>
rect -2162 -1598 2162 1598
<< psubdiff >>
rect -2126 1528 -2030 1562
rect 2030 1528 2126 1562
rect -2126 1466 -2092 1528
rect 2092 1466 2126 1528
rect -2126 -1528 -2092 -1466
rect 2092 -1528 2126 -1466
rect -2126 -1562 -2030 -1528
rect 2030 -1562 2126 -1528
<< psubdiffcont >>
rect -2030 1528 2030 1562
rect -2126 -1466 -2092 1466
rect 2092 -1466 2126 1466
rect -2030 -1562 2030 -1528
<< xpolycontact >>
rect -1996 1000 -1714 1432
rect -1996 -1432 -1714 -1000
rect -1466 1000 -1184 1432
rect -1466 -1432 -1184 -1000
rect -936 1000 -654 1432
rect -936 -1432 -654 -1000
rect -406 1000 -124 1432
rect -406 -1432 -124 -1000
rect 124 1000 406 1432
rect 124 -1432 406 -1000
rect 654 1000 936 1432
rect 654 -1432 936 -1000
rect 1184 1000 1466 1432
rect 1184 -1432 1466 -1000
rect 1714 1000 1996 1432
rect 1714 -1432 1996 -1000
<< xpolyres >>
rect -1996 -1000 -1714 1000
rect -1466 -1000 -1184 1000
rect -936 -1000 -654 1000
rect -406 -1000 -124 1000
rect 124 -1000 406 1000
rect 654 -1000 936 1000
rect 1184 -1000 1466 1000
rect 1714 -1000 1996 1000
<< locali >>
rect -2126 1528 -2030 1562
rect 2030 1528 2126 1562
rect -2126 1466 -2092 1528
rect 2092 1466 2126 1528
rect -2126 -1528 -2092 -1466
rect 2092 -1528 2126 -1466
rect -2126 -1562 -2030 -1528
rect 2030 -1562 2126 -1528
<< viali >>
rect -1980 1017 -1730 1414
rect -1450 1017 -1200 1414
rect -920 1017 -670 1414
rect -390 1017 -140 1414
rect 140 1017 390 1414
rect 670 1017 920 1414
rect 1200 1017 1450 1414
rect 1730 1017 1980 1414
rect -1980 -1414 -1730 -1017
rect -1450 -1414 -1200 -1017
rect -920 -1414 -670 -1017
rect -390 -1414 -140 -1017
rect 140 -1414 390 -1017
rect 670 -1414 920 -1017
rect 1200 -1414 1450 -1017
rect 1730 -1414 1980 -1017
<< metal1 >>
rect -1986 1414 -1724 1426
rect -1986 1017 -1980 1414
rect -1730 1017 -1724 1414
rect -1986 1005 -1724 1017
rect -1456 1414 -1194 1426
rect -1456 1017 -1450 1414
rect -1200 1017 -1194 1414
rect -1456 1005 -1194 1017
rect -926 1414 -664 1426
rect -926 1017 -920 1414
rect -670 1017 -664 1414
rect -926 1005 -664 1017
rect -396 1414 -134 1426
rect -396 1017 -390 1414
rect -140 1017 -134 1414
rect -396 1005 -134 1017
rect 134 1414 396 1426
rect 134 1017 140 1414
rect 390 1017 396 1414
rect 134 1005 396 1017
rect 664 1414 926 1426
rect 664 1017 670 1414
rect 920 1017 926 1414
rect 664 1005 926 1017
rect 1194 1414 1456 1426
rect 1194 1017 1200 1414
rect 1450 1017 1456 1414
rect 1194 1005 1456 1017
rect 1724 1414 1986 1426
rect 1724 1017 1730 1414
rect 1980 1017 1986 1414
rect 1724 1005 1986 1017
rect -1986 -1017 -1724 -1005
rect -1986 -1414 -1980 -1017
rect -1730 -1414 -1724 -1017
rect -1986 -1426 -1724 -1414
rect -1456 -1017 -1194 -1005
rect -1456 -1414 -1450 -1017
rect -1200 -1414 -1194 -1017
rect -1456 -1426 -1194 -1414
rect -926 -1017 -664 -1005
rect -926 -1414 -920 -1017
rect -670 -1414 -664 -1017
rect -926 -1426 -664 -1414
rect -396 -1017 -134 -1005
rect -396 -1414 -390 -1017
rect -140 -1414 -134 -1017
rect -396 -1426 -134 -1414
rect 134 -1017 396 -1005
rect 134 -1414 140 -1017
rect 390 -1414 396 -1017
rect 134 -1426 396 -1414
rect 664 -1017 926 -1005
rect 664 -1414 670 -1017
rect 920 -1414 926 -1017
rect 664 -1426 926 -1414
rect 1194 -1017 1456 -1005
rect 1194 -1414 1200 -1017
rect 1450 -1414 1456 -1017
rect 1194 -1426 1456 -1414
rect 1724 -1017 1986 -1005
rect 1724 -1414 1730 -1017
rect 1980 -1414 1986 -1017
rect 1724 -1426 1986 -1414
<< res1p41 >>
rect -1998 -1002 -1712 1002
rect -1468 -1002 -1182 1002
rect -938 -1002 -652 1002
rect -408 -1002 -122 1002
rect 122 -1002 408 1002
rect 652 -1002 938 1002
rect 1182 -1002 1468 1002
rect 1712 -1002 1998 1002
<< properties >>
string FIXED_BBOX -2109 -1545 2109 1545
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 10 m 1 nx 8 wmin 1.410 lmin 0.50 rho 2000 val 14.451k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
