magic
tech sky130A
magscale 1 2
timestamp 1645462850
<< error_p >>
rect -1996 52 -1714 196
rect -1466 52 -1184 196
rect -936 52 -654 196
rect -406 52 -124 196
rect 124 52 406 196
rect 654 52 936 196
rect 1184 52 1466 196
rect 1714 52 1996 196
<< pwell >>
rect -2162 -3082 2162 3082
<< psubdiff >>
rect -2126 3012 -2030 3046
rect 2030 3012 2126 3046
rect -2126 2950 -2092 3012
rect 2092 2950 2126 3012
rect -2126 -3012 -2092 -2950
rect 2092 -3012 2126 -2950
rect -2126 -3046 -2030 -3012
rect 2030 -3046 2126 -3012
<< psubdiffcont >>
rect -2030 3012 2030 3046
rect -2126 -2950 -2092 2950
rect 2092 -2950 2126 2950
rect -2030 -3046 2030 -3012
<< xpolycontact >>
rect -1996 2484 -1714 2916
rect -1996 52 -1714 484
rect -1466 2484 -1184 2916
rect -1466 52 -1184 484
rect -936 2484 -654 2916
rect -936 52 -654 484
rect -406 2484 -124 2916
rect -406 52 -124 484
rect 124 2484 406 2916
rect 124 52 406 484
rect 654 2484 936 2916
rect 654 52 936 484
rect 1184 2484 1466 2916
rect 1184 52 1466 484
rect 1714 2484 1996 2916
rect 1714 52 1996 484
rect -1996 -484 -1714 -52
rect -1996 -2916 -1714 -2484
rect -1466 -484 -1184 -52
rect -1466 -2916 -1184 -2484
rect -936 -484 -654 -52
rect -936 -2916 -654 -2484
rect -406 -484 -124 -52
rect -406 -2916 -124 -2484
rect 124 -484 406 -52
rect 124 -2916 406 -2484
rect 654 -484 936 -52
rect 654 -2916 936 -2484
rect 1184 -484 1466 -52
rect 1184 -2916 1466 -2484
rect 1714 -484 1996 -52
rect 1714 -2916 1996 -2484
<< xpolyres >>
rect -1996 484 -1714 2484
rect -1466 484 -1184 2484
rect -936 484 -654 2484
rect -406 484 -124 2484
rect 124 484 406 2484
rect 654 484 936 2484
rect 1184 484 1466 2484
rect 1714 484 1996 2484
rect -1996 -2484 -1714 -484
rect -1466 -2484 -1184 -484
rect -936 -2484 -654 -484
rect -406 -2484 -124 -484
rect 124 -2484 406 -484
rect 654 -2484 936 -484
rect 1184 -2484 1466 -484
rect 1714 -2484 1996 -484
<< locali >>
rect -2126 3012 -2030 3046
rect 2030 3012 2126 3046
rect -2126 2950 -2092 3012
rect 2092 2950 2126 3012
rect -2126 -3012 -2092 -2950
rect 2092 -3012 2126 -2950
rect -2126 -3046 -2030 -3012
rect 2030 -3046 2126 -3012
<< viali >>
rect -1980 2501 -1730 2898
rect -1450 2501 -1200 2898
rect -920 2501 -670 2898
rect -390 2501 -140 2898
rect 140 2501 390 2898
rect 670 2501 920 2898
rect 1200 2501 1450 2898
rect 1730 2501 1980 2898
rect -1980 70 -1730 467
rect -1450 70 -1200 467
rect -920 70 -670 467
rect -390 70 -140 467
rect 140 70 390 467
rect 670 70 920 467
rect 1200 70 1450 467
rect 1730 70 1980 467
rect -1980 -467 -1730 -70
rect -1450 -467 -1200 -70
rect -920 -467 -670 -70
rect -390 -467 -140 -70
rect 140 -467 390 -70
rect 670 -467 920 -70
rect 1200 -467 1450 -70
rect 1730 -467 1980 -70
rect -1980 -2898 -1730 -2501
rect -1450 -2898 -1200 -2501
rect -920 -2898 -670 -2501
rect -390 -2898 -140 -2501
rect 140 -2898 390 -2501
rect 670 -2898 920 -2501
rect 1200 -2898 1450 -2501
rect 1730 -2898 1980 -2501
<< metal1 >>
rect -1986 2898 -1724 2910
rect -1986 2501 -1980 2898
rect -1730 2501 -1724 2898
rect -1986 2489 -1724 2501
rect -1456 2898 -1194 2910
rect -1456 2501 -1450 2898
rect -1200 2501 -1194 2898
rect -1456 2489 -1194 2501
rect -926 2898 -664 2910
rect -926 2501 -920 2898
rect -670 2501 -664 2898
rect -926 2489 -664 2501
rect -396 2898 -134 2910
rect -396 2501 -390 2898
rect -140 2501 -134 2898
rect -396 2489 -134 2501
rect 134 2898 396 2910
rect 134 2501 140 2898
rect 390 2501 396 2898
rect 134 2489 396 2501
rect 664 2898 926 2910
rect 664 2501 670 2898
rect 920 2501 926 2898
rect 664 2489 926 2501
rect 1194 2898 1456 2910
rect 1194 2501 1200 2898
rect 1450 2501 1456 2898
rect 1194 2489 1456 2501
rect 1724 2898 1986 2910
rect 1724 2501 1730 2898
rect 1980 2501 1986 2898
rect 1724 2489 1986 2501
rect -1986 467 -1724 479
rect -1986 70 -1980 467
rect -1730 70 -1724 467
rect -1986 58 -1724 70
rect -1456 467 -1194 479
rect -1456 70 -1450 467
rect -1200 70 -1194 467
rect -1456 58 -1194 70
rect -926 467 -664 479
rect -926 70 -920 467
rect -670 70 -664 467
rect -926 58 -664 70
rect -396 467 -134 479
rect -396 70 -390 467
rect -140 70 -134 467
rect -396 58 -134 70
rect 134 467 396 479
rect 134 70 140 467
rect 390 70 396 467
rect 134 58 396 70
rect 664 467 926 479
rect 664 70 670 467
rect 920 70 926 467
rect 664 58 926 70
rect 1194 467 1456 479
rect 1194 70 1200 467
rect 1450 70 1456 467
rect 1194 58 1456 70
rect 1724 467 1986 479
rect 1724 70 1730 467
rect 1980 70 1986 467
rect 1724 58 1986 70
rect -1986 -70 -1724 -58
rect -1986 -467 -1980 -70
rect -1730 -467 -1724 -70
rect -1986 -479 -1724 -467
rect -1456 -70 -1194 -58
rect -1456 -467 -1450 -70
rect -1200 -467 -1194 -70
rect -1456 -479 -1194 -467
rect -926 -70 -664 -58
rect -926 -467 -920 -70
rect -670 -467 -664 -70
rect -926 -479 -664 -467
rect -396 -70 -134 -58
rect -396 -467 -390 -70
rect -140 -467 -134 -70
rect -396 -479 -134 -467
rect 134 -70 396 -58
rect 134 -467 140 -70
rect 390 -467 396 -70
rect 134 -479 396 -467
rect 664 -70 926 -58
rect 664 -467 670 -70
rect 920 -467 926 -70
rect 664 -479 926 -467
rect 1194 -70 1456 -58
rect 1194 -467 1200 -70
rect 1450 -467 1456 -70
rect 1194 -479 1456 -467
rect 1724 -70 1986 -58
rect 1724 -467 1730 -70
rect 1980 -467 1986 -70
rect 1724 -479 1986 -467
rect -1986 -2501 -1724 -2489
rect -1986 -2898 -1980 -2501
rect -1730 -2898 -1724 -2501
rect -1986 -2910 -1724 -2898
rect -1456 -2501 -1194 -2489
rect -1456 -2898 -1450 -2501
rect -1200 -2898 -1194 -2501
rect -1456 -2910 -1194 -2898
rect -926 -2501 -664 -2489
rect -926 -2898 -920 -2501
rect -670 -2898 -664 -2501
rect -926 -2910 -664 -2898
rect -396 -2501 -134 -2489
rect -396 -2898 -390 -2501
rect -140 -2898 -134 -2501
rect -396 -2910 -134 -2898
rect 134 -2501 396 -2489
rect 134 -2898 140 -2501
rect 390 -2898 396 -2501
rect 134 -2910 396 -2898
rect 664 -2501 926 -2489
rect 664 -2898 670 -2501
rect 920 -2898 926 -2501
rect 664 -2910 926 -2898
rect 1194 -2501 1456 -2489
rect 1194 -2898 1200 -2501
rect 1450 -2898 1456 -2501
rect 1194 -2910 1456 -2898
rect 1724 -2501 1986 -2489
rect 1724 -2898 1730 -2501
rect 1980 -2898 1986 -2501
rect 1724 -2910 1986 -2898
<< res1p41 >>
rect -1998 482 -1712 2486
rect -1468 482 -1182 2486
rect -938 482 -652 2486
rect -408 482 -122 2486
rect 122 482 408 2486
rect 652 482 938 2486
rect 1182 482 1468 2486
rect 1712 482 1998 2486
rect -1998 -2486 -1712 -482
rect -1468 -2486 -1182 -482
rect -938 -2486 -652 -482
rect -408 -2486 -122 -482
rect 122 -2486 408 -482
rect 652 -2486 938 -482
rect 1182 -2486 1468 -482
rect 1712 -2486 1998 -482
<< properties >>
string FIXED_BBOX -2109 -3029 2109 3029
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 10 m 2 nx 8 wmin 1.410 lmin 0.50 rho 2000 val 14.451k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
