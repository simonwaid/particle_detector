magic
tech sky130A
timestamp 1646653136
<< pwell >>
rect -1316 -119 1316 119
<< psubdiff >>
rect -1298 84 -1250 101
rect -1144 84 -1096 101
rect -1298 53 -1281 84
rect -1113 53 -1096 84
rect -1298 -84 -1281 -53
rect -1113 -84 -1096 -53
rect -1298 -101 -1250 -84
rect -1144 -101 -1096 -84
rect -1032 84 -984 101
rect -878 84 -830 101
rect -1032 53 -1015 84
rect -847 53 -830 84
rect -1032 -84 -1015 -53
rect -847 -84 -830 -53
rect -1032 -101 -984 -84
rect -878 -101 -830 -84
rect -766 84 -718 101
rect -612 84 -564 101
rect -766 53 -749 84
rect -581 53 -564 84
rect -766 -84 -749 -53
rect -581 -84 -564 -53
rect -766 -101 -718 -84
rect -612 -101 -564 -84
rect -500 84 -452 101
rect -346 84 -298 101
rect -500 53 -483 84
rect -315 53 -298 84
rect -500 -84 -483 -53
rect -315 -84 -298 -53
rect -500 -101 -452 -84
rect -346 -101 -298 -84
rect -234 84 -186 101
rect -80 84 -32 101
rect -234 53 -217 84
rect -49 53 -32 84
rect -234 -84 -217 -53
rect -49 -84 -32 -53
rect -234 -101 -186 -84
rect -80 -101 -32 -84
rect 32 84 80 101
rect 186 84 234 101
rect 32 53 49 84
rect 217 53 234 84
rect 32 -84 49 -53
rect 217 -84 234 -53
rect 32 -101 80 -84
rect 186 -101 234 -84
rect 298 84 346 101
rect 452 84 500 101
rect 298 53 315 84
rect 483 53 500 84
rect 298 -84 315 -53
rect 483 -84 500 -53
rect 298 -101 346 -84
rect 452 -101 500 -84
rect 564 84 612 101
rect 718 84 766 101
rect 564 53 581 84
rect 749 53 766 84
rect 564 -84 581 -53
rect 749 -84 766 -53
rect 564 -101 612 -84
rect 718 -101 766 -84
rect 830 84 878 101
rect 984 84 1032 101
rect 830 53 847 84
rect 1015 53 1032 84
rect 830 -84 847 -53
rect 1015 -84 1032 -53
rect 830 -101 878 -84
rect 984 -101 1032 -84
rect 1096 84 1144 101
rect 1250 84 1298 101
rect 1096 53 1113 84
rect 1281 53 1298 84
rect 1096 -84 1113 -53
rect 1281 -84 1298 -53
rect 1096 -101 1144 -84
rect 1250 -101 1298 -84
<< psubdiffcont >>
rect -1250 84 -1144 101
rect -1298 -53 -1281 53
rect -1113 -53 -1096 53
rect -1250 -101 -1144 -84
rect -984 84 -878 101
rect -1032 -53 -1015 53
rect -847 -53 -830 53
rect -984 -101 -878 -84
rect -718 84 -612 101
rect -766 -53 -749 53
rect -581 -53 -564 53
rect -718 -101 -612 -84
rect -452 84 -346 101
rect -500 -53 -483 53
rect -315 -53 -298 53
rect -452 -101 -346 -84
rect -186 84 -80 101
rect -234 -53 -217 53
rect -49 -53 -32 53
rect -186 -101 -80 -84
rect 80 84 186 101
rect 32 -53 49 53
rect 217 -53 234 53
rect 80 -101 186 -84
rect 346 84 452 101
rect 298 -53 315 53
rect 483 -53 500 53
rect 346 -101 452 -84
rect 612 84 718 101
rect 564 -53 581 53
rect 749 -53 766 53
rect 612 -101 718 -84
rect 878 84 984 101
rect 830 -53 847 53
rect 1015 -53 1032 53
rect 878 -101 984 -84
rect 1144 84 1250 101
rect 1096 -53 1113 53
rect 1281 -53 1298 53
rect 1144 -101 1250 -84
<< ndiode >>
rect -1247 44 -1147 50
rect -1247 -44 -1241 44
rect -1153 -44 -1147 44
rect -1247 -50 -1147 -44
rect -981 44 -881 50
rect -981 -44 -975 44
rect -887 -44 -881 44
rect -981 -50 -881 -44
rect -715 44 -615 50
rect -715 -44 -709 44
rect -621 -44 -615 44
rect -715 -50 -615 -44
rect -449 44 -349 50
rect -449 -44 -443 44
rect -355 -44 -349 44
rect -449 -50 -349 -44
rect -183 44 -83 50
rect -183 -44 -177 44
rect -89 -44 -83 44
rect -183 -50 -83 -44
rect 83 44 183 50
rect 83 -44 89 44
rect 177 -44 183 44
rect 83 -50 183 -44
rect 349 44 449 50
rect 349 -44 355 44
rect 443 -44 449 44
rect 349 -50 449 -44
rect 615 44 715 50
rect 615 -44 621 44
rect 709 -44 715 44
rect 615 -50 715 -44
rect 881 44 981 50
rect 881 -44 887 44
rect 975 -44 981 44
rect 881 -50 981 -44
rect 1147 44 1247 50
rect 1147 -44 1153 44
rect 1241 -44 1247 44
rect 1147 -50 1247 -44
<< ndiodec >>
rect -1241 -44 -1153 44
rect -975 -44 -887 44
rect -709 -44 -621 44
rect -443 -44 -355 44
rect -177 -44 -89 44
rect 89 -44 177 44
rect 355 -44 443 44
rect 621 -44 709 44
rect 887 -44 975 44
rect 1153 -44 1241 44
<< locali >>
rect -1298 84 -1250 101
rect -1144 84 -1096 101
rect -1298 53 -1281 84
rect -1113 53 -1096 84
rect -1249 -44 -1241 44
rect -1153 -44 -1145 44
rect -1298 -84 -1281 -53
rect -1113 -84 -1096 -53
rect -1298 -101 -1250 -84
rect -1144 -101 -1096 -84
rect -1032 84 -984 101
rect -878 84 -830 101
rect -1032 53 -1015 84
rect -847 53 -830 84
rect -983 -44 -975 44
rect -887 -44 -879 44
rect -1032 -84 -1015 -53
rect -847 -84 -830 -53
rect -1032 -101 -984 -84
rect -878 -101 -830 -84
rect -766 84 -718 101
rect -612 84 -564 101
rect -766 53 -749 84
rect -581 53 -564 84
rect -717 -44 -709 44
rect -621 -44 -613 44
rect -766 -84 -749 -53
rect -581 -84 -564 -53
rect -766 -101 -718 -84
rect -612 -101 -564 -84
rect -500 84 -452 101
rect -346 84 -298 101
rect -500 53 -483 84
rect -315 53 -298 84
rect -451 -44 -443 44
rect -355 -44 -347 44
rect -500 -84 -483 -53
rect -315 -84 -298 -53
rect -500 -101 -452 -84
rect -346 -101 -298 -84
rect -234 84 -186 101
rect -80 84 -32 101
rect -234 53 -217 84
rect -49 53 -32 84
rect -185 -44 -177 44
rect -89 -44 -81 44
rect -234 -84 -217 -53
rect -49 -84 -32 -53
rect -234 -101 -186 -84
rect -80 -101 -32 -84
rect 32 84 80 101
rect 186 84 234 101
rect 32 53 49 84
rect 217 53 234 84
rect 81 -44 89 44
rect 177 -44 185 44
rect 32 -84 49 -53
rect 217 -84 234 -53
rect 32 -101 80 -84
rect 186 -101 234 -84
rect 298 84 346 101
rect 452 84 500 101
rect 298 53 315 84
rect 483 53 500 84
rect 347 -44 355 44
rect 443 -44 451 44
rect 298 -84 315 -53
rect 483 -84 500 -53
rect 298 -101 346 -84
rect 452 -101 500 -84
rect 564 84 612 101
rect 718 84 766 101
rect 564 53 581 84
rect 749 53 766 84
rect 613 -44 621 44
rect 709 -44 717 44
rect 564 -84 581 -53
rect 749 -84 766 -53
rect 564 -101 612 -84
rect 718 -101 766 -84
rect 830 84 878 101
rect 984 84 1032 101
rect 830 53 847 84
rect 1015 53 1032 84
rect 879 -44 887 44
rect 975 -44 983 44
rect 830 -84 847 -53
rect 1015 -84 1032 -53
rect 830 -101 878 -84
rect 984 -101 1032 -84
rect 1096 84 1144 101
rect 1250 84 1298 101
rect 1096 53 1113 84
rect 1281 53 1298 84
rect 1145 -44 1153 44
rect 1241 -44 1249 44
rect 1096 -84 1113 -53
rect 1281 -84 1298 -53
rect 1096 -101 1144 -84
rect 1250 -101 1298 -84
<< viali >>
rect -1241 -44 -1153 44
rect -975 -44 -887 44
rect -709 -44 -621 44
rect -443 -44 -355 44
rect -177 -44 -89 44
rect 89 -44 177 44
rect 355 -44 443 44
rect 621 -44 709 44
rect 887 -44 975 44
rect 1153 -44 1241 44
<< metal1 >>
rect -1247 44 -1147 47
rect -1247 -44 -1241 44
rect -1153 -44 -1147 44
rect -1247 -47 -1147 -44
rect -981 44 -881 47
rect -981 -44 -975 44
rect -887 -44 -881 44
rect -981 -47 -881 -44
rect -715 44 -615 47
rect -715 -44 -709 44
rect -621 -44 -615 44
rect -715 -47 -615 -44
rect -449 44 -349 47
rect -449 -44 -443 44
rect -355 -44 -349 44
rect -449 -47 -349 -44
rect -183 44 -83 47
rect -183 -44 -177 44
rect -89 -44 -83 44
rect -183 -47 -83 -44
rect 83 44 183 47
rect 83 -44 89 44
rect 177 -44 183 44
rect 83 -47 183 -44
rect 349 44 449 47
rect 349 -44 355 44
rect 443 -44 449 44
rect 349 -47 449 -44
rect 615 44 715 47
rect 615 -44 621 44
rect 709 -44 715 44
rect 615 -47 715 -44
rect 881 44 981 47
rect 881 -44 887 44
rect 975 -44 981 44
rect 881 -47 981 -44
rect 1147 44 1247 47
rect 1147 -44 1153 44
rect 1241 -44 1247 44
rect 1147 -47 1247 -44
<< properties >>
string FIXED_BBOX 1104 -92 1289 92
string gencell sky130_fd_pr__diode_pw2nd_05v5
string library sky130
string parameters w 1 l 1 area 1.0 peri 4.0 nx 10 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
