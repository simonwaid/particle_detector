magic
tech sky130A
magscale 1 2
timestamp 1647868710
<< pwell >>
rect -19838 7542 -19676 7608
rect -19838 7032 -19676 7098
<< poly >>
rect -19838 7592 -19676 7608
rect -19838 7558 -19822 7592
rect -19788 7558 -19676 7592
rect -19838 7542 -19676 7558
rect -19838 7082 -19676 7098
rect -19838 7048 -19726 7082
rect -19692 7048 -19676 7082
rect -19838 7032 -19676 7048
<< polycont >>
rect -19822 7558 -19788 7592
rect -19726 7048 -19692 7082
<< locali >>
rect -19838 7558 -19822 7592
rect -19788 7558 -19676 7592
rect -19838 7048 -19726 7082
rect -19692 7048 -19676 7082
rect -19540 6960 -19470 7690
rect -20100 6860 -19470 6960
rect -19540 5510 -19470 6860
<< viali >>
rect -19822 7558 -19788 7592
rect -19726 7048 -19692 7082
<< metal1 >>
rect -21110 13500 -21100 15200
rect -14440 13500 -14430 15200
rect -19850 7550 -19840 7710
rect -19680 7630 -19670 7710
rect -19680 7550 -19470 7630
rect -19780 7520 -19734 7550
rect -19890 7120 -19880 7280
rect -19826 7120 -19816 7280
rect -19698 7120 -19688 7280
rect -19634 7120 -19624 7280
rect -19780 7090 -19734 7120
rect -19950 7082 -19460 7090
rect -19950 7048 -19726 7082
rect -19692 7048 -19460 7082
rect -19950 6730 -19460 7048
rect -19852 6538 -19842 6698
rect -19788 6538 -19778 6698
rect -16680 6460 -14280 6840
rect -20010 6298 -20000 6458
rect -19946 6298 -19936 6458
rect -19694 6298 -19684 6458
rect -19630 6298 -19620 6458
rect -19950 6110 -19470 6270
rect -20010 5920 -20000 6080
rect -19946 5920 -19936 6080
rect -19694 5920 -19684 6080
rect -19630 5920 -19620 6080
rect -19852 5680 -19842 5840
rect -19788 5680 -19778 5840
rect -19950 5570 -19470 5650
rect -120 1040 40 6040
<< via1 >>
rect -21100 13500 -14440 15200
rect -19840 7592 -19680 7710
rect -19840 7558 -19822 7592
rect -19822 7558 -19788 7592
rect -19788 7558 -19680 7592
rect -19840 7550 -19680 7558
rect -19880 7120 -19826 7280
rect -19688 7120 -19634 7280
rect -19842 6538 -19788 6698
rect -20000 6298 -19946 6458
rect -19684 6298 -19630 6458
rect -20000 5920 -19946 6080
rect -19684 5920 -19630 6080
rect -19842 5680 -19788 5840
<< metal2 >>
rect -21100 15200 -14440 15210
rect -21100 13490 -14440 13500
rect -300 13460 60 13470
rect -1160 12780 -800 12790
rect -15460 11640 -15100 11660
rect -21080 11310 -20960 11420
rect -15460 11280 -15440 11640
rect -15120 11280 -15100 11640
rect -21150 10590 -20890 10600
rect -21150 10290 -20890 10300
rect -21090 9740 -20940 10290
rect -15460 9300 -15100 11280
rect -14760 10580 -14400 12280
rect -14760 10400 -14280 10580
rect -1160 9300 -800 12420
rect -300 10760 60 13100
rect -300 10400 54680 10760
rect -15460 9120 -14280 9300
rect -1160 8940 54700 9300
rect -20220 7920 -19680 7930
rect -20220 7780 -19830 7920
rect -19690 7780 -19680 7920
rect -20220 7770 -19680 7780
rect -19840 7710 -19680 7770
rect -19840 7540 -19680 7550
rect -19900 7280 -19630 7290
rect -19900 7120 -19880 7280
rect -19826 7120 -19688 7280
rect -19634 7120 -19630 7280
rect -19900 7110 -19630 7120
rect -19900 6750 -19720 7110
rect -19900 6698 -19730 6750
rect -19900 6538 -19842 6698
rect -19788 6538 -19730 6698
rect -20100 6458 -19940 6470
rect -20100 6298 -20000 6458
rect -19946 6298 -19940 6458
rect -20100 6080 -19940 6298
rect -20100 5920 -20000 6080
rect -19946 5920 -19940 6080
rect -20100 5520 -19940 5920
rect -19900 5840 -19730 6538
rect -19900 5680 -19842 5840
rect -19788 5680 -19730 5840
rect -19900 5670 -19730 5680
rect -19690 6458 -19530 6470
rect -19690 6298 -19684 6458
rect -19630 6298 -19530 6458
rect -19690 6080 -19530 6298
rect -19690 5920 -19684 6080
rect -19630 5920 -19530 6080
rect -19690 5840 -19530 5920
rect -19690 5520 -19340 5840
rect -20100 5360 -19340 5520
rect -19570 5300 -19340 5360
<< via2 >>
rect -21100 13500 -14440 15200
rect -300 13100 60 13460
rect -1160 12420 -800 12780
rect -15440 11280 -15120 11640
rect -21150 10300 -20890 10590
rect -19830 7780 -19690 7920
<< metal3 >>
rect -21110 15200 -14430 15205
rect -21110 13500 -21100 15200
rect -14440 13500 -14430 15200
rect -13930 14260 -13920 14960
rect -2520 14260 -2510 14960
rect 390 14260 400 14960
rect 11800 14260 11810 14960
rect 14650 14260 14660 14960
rect 26060 14260 26070 14960
rect 28890 14260 28900 14960
rect 40300 14260 40310 14960
rect 43150 14260 43160 14960
rect 54560 14260 54570 14960
rect -21110 13495 -14430 13500
rect -310 13460 70 13465
rect -310 13100 -300 13460
rect 60 13100 70 13460
rect -310 13095 70 13100
rect -1170 12780 -790 12785
rect -1170 12420 -1160 12780
rect -800 12420 -790 12780
rect -1170 12415 -790 12420
rect -15450 11640 -15110 11645
rect -15450 11280 -15440 11640
rect -15120 11280 -15110 11640
rect -15450 11275 -15110 11280
rect -26280 10780 -25380 11120
rect -21610 10780 -19680 10910
rect -21160 10590 -20880 10595
rect -21160 10300 -21150 10590
rect -20890 10300 -20880 10590
rect -21160 10295 -20880 10300
rect -19840 7920 -19680 10780
rect -12280 8500 -12000 8690
rect 2030 8460 2280 8660
rect -19840 7780 -19830 7920
rect -19690 7780 -19680 7920
rect -19840 7770 -19680 7780
rect -18488 1660 -17582 2134
rect -19490 440 -19480 1660
rect -16640 440 -16630 1660
rect -14310 20 -14300 960
rect 56940 20 56950 960
<< via3 >>
rect -21100 13500 -14440 15200
rect -13920 14260 -2520 14960
rect 400 14260 11800 14960
rect 14660 14260 26060 14960
rect 28900 14260 40300 14960
rect 43160 14260 54560 14960
rect -300 13100 60 13460
rect -1160 12420 -800 12780
rect -15440 11280 -15120 11640
rect -21150 10300 -20890 10590
rect -19480 440 -16640 1660
rect -14300 20 56940 960
<< metal4 >>
rect -21101 15200 -14439 15201
rect -21101 13500 -21100 15200
rect -14440 13500 -14439 15200
rect -13921 14960 -2519 14961
rect -13921 14260 -13920 14960
rect -2520 14260 -2519 14960
rect -13921 14259 -2519 14260
rect 399 14960 11801 14961
rect 399 14260 400 14960
rect 11800 14260 11801 14960
rect 399 14259 11801 14260
rect 14659 14960 26061 14961
rect 14659 14260 14660 14960
rect 26060 14260 26061 14960
rect 14659 14259 26061 14260
rect 28899 14960 40301 14961
rect 28899 14260 28900 14960
rect 40300 14260 40301 14960
rect 28899 14259 40301 14260
rect 43159 14960 54561 14961
rect 43159 14260 43160 14960
rect 54560 14260 54561 14960
rect 43159 14259 54561 14260
rect -21101 13499 -14439 13500
rect -301 13460 61 13461
rect -2360 13100 -300 13460
rect 60 13100 61 13460
rect -2360 12900 -2340 13100
rect -301 13099 61 13100
rect -300 13080 60 13099
rect 54740 12900 55850 13460
rect -1161 12780 -799 12781
rect -2360 12420 -1160 12780
rect -800 12420 -799 12780
rect -2360 12220 -2320 12420
rect -1161 12419 -799 12420
rect -1160 12400 -800 12419
rect 54740 12220 55850 12780
rect -15441 11640 -15119 11641
rect -15441 11280 -15440 11640
rect -15120 11280 -15119 11640
rect -15441 11279 -15119 11280
rect -30140 10200 -21350 10760
rect -21151 10590 -20889 10591
rect -21151 10300 -21150 10590
rect -20890 10300 -20889 10590
rect -21151 10299 -20889 10300
rect -30140 10100 -20900 10200
rect -19481 1660 -16639 1661
rect -19481 440 -19480 1660
rect -16640 440 -16639 1660
rect -19481 439 -16639 440
rect -14301 960 56941 961
rect -14301 20 -14300 960
rect 56940 20 56941 960
rect -14301 19 56941 20
<< via4 >>
rect -21100 13500 -14440 15200
rect -13920 14260 -2520 14960
rect 400 14260 11800 14960
rect 14660 14260 26060 14960
rect 28900 14260 40300 14960
rect 43160 14260 54560 14960
rect -21150 10300 -20890 10590
rect -19480 440 -16640 1660
rect -14300 20 56940 960
<< metal5 >>
rect -21124 15220 -14416 15224
rect -30160 15200 57000 15220
rect -30160 13500 -21100 15200
rect -14440 14960 57000 15200
rect -14440 14260 -13920 14960
rect -2520 14260 400 14960
rect 11800 14260 14660 14960
rect 26060 14260 28900 14960
rect 40300 14260 43160 14960
rect 54560 14260 57000 14960
rect -14440 13500 57000 14260
rect -30160 12500 57000 13500
rect -21180 10590 -20850 10620
rect -21180 10300 -21150 10590
rect -20890 10300 -20850 10590
rect -21180 9980 -20850 10300
rect -13920 9980 -12900 12500
rect -6820 10000 -5800 12500
rect 580 10020 1600 12500
rect 8100 9940 9120 12500
rect 15640 9920 16660 12500
rect 23420 9980 24440 12500
rect 31200 9980 32220 12500
rect 40060 10040 41080 12500
rect 49480 10000 50500 12500
rect -22620 9330 -21510 9720
rect -28540 2660 -15540 3640
rect -14000 2660 -12980 4920
rect -6580 2660 -5560 4920
rect 780 2660 1800 5060
rect 8520 2660 9540 5160
rect 16060 2660 17080 5180
rect 24000 2660 25020 5060
rect 31660 2660 32680 5300
rect 40040 2660 41060 4880
rect 48700 2660 49720 4840
rect -29980 1660 57040 2660
rect -29980 440 -19480 1660
rect -16640 960 57040 1660
rect -16640 440 -14300 960
rect -29980 20 -14300 440
rect 56940 20 57040 960
rect -29980 -60 57040 20
use outd_stage1  outd_stage1_0
timestamp 1647868710
transform 1 0 -19480 0 1 1680
box -1660 -880 5040 12406
use outd_stage2  outd_stage2_0
timestamp 1647868710
transform 1 0 -14290 0 1 880
box -30 -880 14232 14120
use outd_stage3  outd_stage3_0
timestamp 1647868710
transform 1 0 20 0 1 20
box -20 -20 56992 14980
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_0
timestamp 1647868710
transform 0 -1 -23680 1 0 12740
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_1
timestamp 1647868710
transform 0 -1 -28120 1 0 12750
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1647868710
transform 0 -1 -11199 1 0 6791
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_1
timestamp 1647868710
transform 0 -1 -3999 1 0 6791
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_2
timestamp 1647868710
transform 0 -1 3421 1 0 6771
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_3
timestamp 1647868710
transform 0 -1 11001 1 0 6751
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_4
timestamp 1647868710
transform 0 -1 18501 1 0 6751
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_5
timestamp 1647868710
transform 0 -1 26261 1 0 6771
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_6
timestamp 1647868710
transform 0 -1 33781 1 0 6771
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_7
timestamp 1647868710
transform 0 -1 42561 1 0 6831
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_8
timestamp 1647868710
transform 0 -1 50901 1 0 6811
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_9
timestamp 1647868710
transform 0 1 -18659 -1 0 6793
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_10
timestamp 1647868710
transform 0 1 -25439 -1 0 6813
box -3351 -3101 3373 3101
use sky130_fd_pr__nfet_01v8_DJG2KN  sky130_fd_pr__nfet_01v8_DJG2KN_0
timestamp 1647868710
transform 1 0 -19815 0 1 6189
box -325 -719 325 719
use sky130_fd_pr__nfet_01v8_LH2JGW  sky130_fd_pr__nfet_01v8_LH2JGW_0
timestamp 1647868710
transform 1 0 -19757 0 1 7320
box -263 -410 263 410
<< labels >>
rlabel metal2 -20210 7780 -20050 7920 1 I_Bias
rlabel metal2 -21080 11310 -20960 11420 1 InputSignal
rlabel metal2 -21080 9750 -20950 9860 1 InputRef
rlabel metal2 -15390 10580 -15190 10730 1 V_da1_P
rlabel metal2 -14690 10610 -14490 10760 1 V_da1_N
rlabel metal5 -29610 520 -28750 1280 1 VN
rlabel metal5 -29780 13450 -28910 14580 1 VP
rlabel metal2 -1090 11190 -910 11400 1 V_da2_P
rlabel metal2 -170 11220 10 11430 1 V_da2_N
rlabel metal4 55470 12270 55650 12440 1 OutputP
rlabel metal4 55470 12940 55650 13140 3 OutputN
rlabel metal3 -12280 8500 -12000 8690 1 VM1_D
rlabel metal3 2030 8460 2280 8660 1 VM14D
<< end >>
