* SPICE3 file created from outd_stage1.ext - technology: sky130A

X0 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 isource_out m1_260_8900# m1_n1500_10180# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 m1_n1500_10180# m1_260_8900# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X39 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X40 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X41 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X42 isource_out m1_1860_8350# m1_1830_10170# isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X43 m1_1830_10170# m1_1860_8350# isource_out isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 m1_n1500_10180# dw_70_8020# VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X45 m1_n1500_10180# dw_70_8020# VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X46 m1_n1500_10180# dw_70_8020# VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X47 m1_n1500_10180# dw_70_8020# VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X48 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X51 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X53 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X56 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X57 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X58 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X59 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X61 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X64 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X65 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X66 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X67 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X69 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X70 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X72 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X75 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X76 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X77 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X80 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X83 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X85 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X90 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X92 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X93 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X94 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X98 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X99 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X100 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X101 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X102 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X104 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X105 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X106 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X107 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X108 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X109 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X110 isource_out outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X111 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X112 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X113 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X114 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X115 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X116 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X117 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X118 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X119 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X120 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X121 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X122 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X123 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X124 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X125 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X126 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X127 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X128 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X129 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X130 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X131 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X132 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X133 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X134 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X135 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X136 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X137 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X138 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X139 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X140 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X141 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X142 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X143 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X145 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X146 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X147 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X148 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X149 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X150 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X151 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X152 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X153 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X154 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X155 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X156 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X157 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X158 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X159 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X160 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X161 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X162 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X163 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X164 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X165 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X166 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X167 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X168 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X169 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X170 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X171 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X172 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X173 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X174 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X175 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X176 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X177 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X178 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X179 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X180 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X181 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X182 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X183 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X184 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X185 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X186 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X187 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X188 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X189 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X190 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X191 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X192 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X193 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X194 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X195 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X196 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X197 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X198 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X199 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X200 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X201 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X202 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X203 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X204 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X205 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X206 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X207 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X208 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X209 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X210 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X211 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X212 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X213 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X214 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X215 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X216 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X217 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X218 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X219 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X220 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X221 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X222 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X223 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X224 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X225 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X226 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X227 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X228 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X229 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X230 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X231 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X232 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X233 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X234 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X235 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X236 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X237 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X238 VN outd_cmirror_64t_0/m1_0_80# outd_cmirror_64t_0/m1_220_5610# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X239 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X240 m1_1830_10170# dw_70_8020# VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X241 m1_1830_10170# dw_70_8020# VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X242 m1_1830_10170# dw_70_8020# VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X243 m1_1830_10170# dw_70_8020# VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
