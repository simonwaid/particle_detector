magic
tech sky130A
magscale 1 2
timestamp 1646234887
<< pwell >>
rect -1431 -1028 1431 1028
<< nmos >>
rect -1235 418 -1135 818
rect -1077 418 -977 818
rect -919 418 -819 818
rect -761 418 -661 818
rect -603 418 -503 818
rect -445 418 -345 818
rect -287 418 -187 818
rect -129 418 -29 818
rect 29 418 129 818
rect 187 418 287 818
rect 345 418 445 818
rect 503 418 603 818
rect 661 418 761 818
rect 819 418 919 818
rect 977 418 1077 818
rect 1135 418 1235 818
rect -1235 -200 -1135 200
rect -1077 -200 -977 200
rect -919 -200 -819 200
rect -761 -200 -661 200
rect -603 -200 -503 200
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
rect 503 -200 603 200
rect 661 -200 761 200
rect 819 -200 919 200
rect 977 -200 1077 200
rect 1135 -200 1235 200
rect -1235 -818 -1135 -418
rect -1077 -818 -977 -418
rect -919 -818 -819 -418
rect -761 -818 -661 -418
rect -603 -818 -503 -418
rect -445 -818 -345 -418
rect -287 -818 -187 -418
rect -129 -818 -29 -418
rect 29 -818 129 -418
rect 187 -818 287 -418
rect 345 -818 445 -418
rect 503 -818 603 -418
rect 661 -818 761 -418
rect 819 -818 919 -418
rect 977 -818 1077 -418
rect 1135 -818 1235 -418
<< ndiff >>
rect -1293 806 -1235 818
rect -1293 430 -1281 806
rect -1247 430 -1235 806
rect -1293 418 -1235 430
rect -1135 806 -1077 818
rect -1135 430 -1123 806
rect -1089 430 -1077 806
rect -1135 418 -1077 430
rect -977 806 -919 818
rect -977 430 -965 806
rect -931 430 -919 806
rect -977 418 -919 430
rect -819 806 -761 818
rect -819 430 -807 806
rect -773 430 -761 806
rect -819 418 -761 430
rect -661 806 -603 818
rect -661 430 -649 806
rect -615 430 -603 806
rect -661 418 -603 430
rect -503 806 -445 818
rect -503 430 -491 806
rect -457 430 -445 806
rect -503 418 -445 430
rect -345 806 -287 818
rect -345 430 -333 806
rect -299 430 -287 806
rect -345 418 -287 430
rect -187 806 -129 818
rect -187 430 -175 806
rect -141 430 -129 806
rect -187 418 -129 430
rect -29 806 29 818
rect -29 430 -17 806
rect 17 430 29 806
rect -29 418 29 430
rect 129 806 187 818
rect 129 430 141 806
rect 175 430 187 806
rect 129 418 187 430
rect 287 806 345 818
rect 287 430 299 806
rect 333 430 345 806
rect 287 418 345 430
rect 445 806 503 818
rect 445 430 457 806
rect 491 430 503 806
rect 445 418 503 430
rect 603 806 661 818
rect 603 430 615 806
rect 649 430 661 806
rect 603 418 661 430
rect 761 806 819 818
rect 761 430 773 806
rect 807 430 819 806
rect 761 418 819 430
rect 919 806 977 818
rect 919 430 931 806
rect 965 430 977 806
rect 919 418 977 430
rect 1077 806 1135 818
rect 1077 430 1089 806
rect 1123 430 1135 806
rect 1077 418 1135 430
rect 1235 806 1293 818
rect 1235 430 1247 806
rect 1281 430 1293 806
rect 1235 418 1293 430
rect -1293 188 -1235 200
rect -1293 -188 -1281 188
rect -1247 -188 -1235 188
rect -1293 -200 -1235 -188
rect -1135 188 -1077 200
rect -1135 -188 -1123 188
rect -1089 -188 -1077 188
rect -1135 -200 -1077 -188
rect -977 188 -919 200
rect -977 -188 -965 188
rect -931 -188 -919 188
rect -977 -200 -919 -188
rect -819 188 -761 200
rect -819 -188 -807 188
rect -773 -188 -761 188
rect -819 -200 -761 -188
rect -661 188 -603 200
rect -661 -188 -649 188
rect -615 -188 -603 188
rect -661 -200 -603 -188
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
rect 603 188 661 200
rect 603 -188 615 188
rect 649 -188 661 188
rect 603 -200 661 -188
rect 761 188 819 200
rect 761 -188 773 188
rect 807 -188 819 188
rect 761 -200 819 -188
rect 919 188 977 200
rect 919 -188 931 188
rect 965 -188 977 188
rect 919 -200 977 -188
rect 1077 188 1135 200
rect 1077 -188 1089 188
rect 1123 -188 1135 188
rect 1077 -200 1135 -188
rect 1235 188 1293 200
rect 1235 -188 1247 188
rect 1281 -188 1293 188
rect 1235 -200 1293 -188
rect -1293 -430 -1235 -418
rect -1293 -806 -1281 -430
rect -1247 -806 -1235 -430
rect -1293 -818 -1235 -806
rect -1135 -430 -1077 -418
rect -1135 -806 -1123 -430
rect -1089 -806 -1077 -430
rect -1135 -818 -1077 -806
rect -977 -430 -919 -418
rect -977 -806 -965 -430
rect -931 -806 -919 -430
rect -977 -818 -919 -806
rect -819 -430 -761 -418
rect -819 -806 -807 -430
rect -773 -806 -761 -430
rect -819 -818 -761 -806
rect -661 -430 -603 -418
rect -661 -806 -649 -430
rect -615 -806 -603 -430
rect -661 -818 -603 -806
rect -503 -430 -445 -418
rect -503 -806 -491 -430
rect -457 -806 -445 -430
rect -503 -818 -445 -806
rect -345 -430 -287 -418
rect -345 -806 -333 -430
rect -299 -806 -287 -430
rect -345 -818 -287 -806
rect -187 -430 -129 -418
rect -187 -806 -175 -430
rect -141 -806 -129 -430
rect -187 -818 -129 -806
rect -29 -430 29 -418
rect -29 -806 -17 -430
rect 17 -806 29 -430
rect -29 -818 29 -806
rect 129 -430 187 -418
rect 129 -806 141 -430
rect 175 -806 187 -430
rect 129 -818 187 -806
rect 287 -430 345 -418
rect 287 -806 299 -430
rect 333 -806 345 -430
rect 287 -818 345 -806
rect 445 -430 503 -418
rect 445 -806 457 -430
rect 491 -806 503 -430
rect 445 -818 503 -806
rect 603 -430 661 -418
rect 603 -806 615 -430
rect 649 -806 661 -430
rect 603 -818 661 -806
rect 761 -430 819 -418
rect 761 -806 773 -430
rect 807 -806 819 -430
rect 761 -818 819 -806
rect 919 -430 977 -418
rect 919 -806 931 -430
rect 965 -806 977 -430
rect 919 -818 977 -806
rect 1077 -430 1135 -418
rect 1077 -806 1089 -430
rect 1123 -806 1135 -430
rect 1077 -818 1135 -806
rect 1235 -430 1293 -418
rect 1235 -806 1247 -430
rect 1281 -806 1293 -430
rect 1235 -818 1293 -806
<< ndiffc >>
rect -1281 430 -1247 806
rect -1123 430 -1089 806
rect -965 430 -931 806
rect -807 430 -773 806
rect -649 430 -615 806
rect -491 430 -457 806
rect -333 430 -299 806
rect -175 430 -141 806
rect -17 430 17 806
rect 141 430 175 806
rect 299 430 333 806
rect 457 430 491 806
rect 615 430 649 806
rect 773 430 807 806
rect 931 430 965 806
rect 1089 430 1123 806
rect 1247 430 1281 806
rect -1281 -188 -1247 188
rect -1123 -188 -1089 188
rect -965 -188 -931 188
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect 931 -188 965 188
rect 1089 -188 1123 188
rect 1247 -188 1281 188
rect -1281 -806 -1247 -430
rect -1123 -806 -1089 -430
rect -965 -806 -931 -430
rect -807 -806 -773 -430
rect -649 -806 -615 -430
rect -491 -806 -457 -430
rect -333 -806 -299 -430
rect -175 -806 -141 -430
rect -17 -806 17 -430
rect 141 -806 175 -430
rect 299 -806 333 -430
rect 457 -806 491 -430
rect 615 -806 649 -430
rect 773 -806 807 -430
rect 931 -806 965 -430
rect 1089 -806 1123 -430
rect 1247 -806 1281 -430
<< psubdiff >>
rect -1395 958 -1299 992
rect 1299 958 1395 992
rect -1395 896 -1361 958
rect 1361 896 1395 958
rect -1395 -958 -1361 -896
rect 1361 -958 1395 -896
rect -1395 -992 -1299 -958
rect 1299 -992 1395 -958
<< psubdiffcont >>
rect -1299 958 1299 992
rect -1395 -896 -1361 896
rect 1361 -896 1395 896
rect -1299 -992 1299 -958
<< poly >>
rect -1235 890 -1135 906
rect -1235 856 -1219 890
rect -1151 856 -1135 890
rect -1235 818 -1135 856
rect -1077 890 -977 906
rect -1077 856 -1061 890
rect -993 856 -977 890
rect -1077 818 -977 856
rect -919 890 -819 906
rect -919 856 -903 890
rect -835 856 -819 890
rect -919 818 -819 856
rect -761 890 -661 906
rect -761 856 -745 890
rect -677 856 -661 890
rect -761 818 -661 856
rect -603 890 -503 906
rect -603 856 -587 890
rect -519 856 -503 890
rect -603 818 -503 856
rect -445 890 -345 906
rect -445 856 -429 890
rect -361 856 -345 890
rect -445 818 -345 856
rect -287 890 -187 906
rect -287 856 -271 890
rect -203 856 -187 890
rect -287 818 -187 856
rect -129 890 -29 906
rect -129 856 -113 890
rect -45 856 -29 890
rect -129 818 -29 856
rect 29 890 129 906
rect 29 856 45 890
rect 113 856 129 890
rect 29 818 129 856
rect 187 890 287 906
rect 187 856 203 890
rect 271 856 287 890
rect 187 818 287 856
rect 345 890 445 906
rect 345 856 361 890
rect 429 856 445 890
rect 345 818 445 856
rect 503 890 603 906
rect 503 856 519 890
rect 587 856 603 890
rect 503 818 603 856
rect 661 890 761 906
rect 661 856 677 890
rect 745 856 761 890
rect 661 818 761 856
rect 819 890 919 906
rect 819 856 835 890
rect 903 856 919 890
rect 819 818 919 856
rect 977 890 1077 906
rect 977 856 993 890
rect 1061 856 1077 890
rect 977 818 1077 856
rect 1135 890 1235 906
rect 1135 856 1151 890
rect 1219 856 1235 890
rect 1135 818 1235 856
rect -1235 380 -1135 418
rect -1235 346 -1219 380
rect -1151 346 -1135 380
rect -1235 330 -1135 346
rect -1077 380 -977 418
rect -1077 346 -1061 380
rect -993 346 -977 380
rect -1077 330 -977 346
rect -919 380 -819 418
rect -919 346 -903 380
rect -835 346 -819 380
rect -919 330 -819 346
rect -761 380 -661 418
rect -761 346 -745 380
rect -677 346 -661 380
rect -761 330 -661 346
rect -603 380 -503 418
rect -603 346 -587 380
rect -519 346 -503 380
rect -603 330 -503 346
rect -445 380 -345 418
rect -445 346 -429 380
rect -361 346 -345 380
rect -445 330 -345 346
rect -287 380 -187 418
rect -287 346 -271 380
rect -203 346 -187 380
rect -287 330 -187 346
rect -129 380 -29 418
rect -129 346 -113 380
rect -45 346 -29 380
rect -129 330 -29 346
rect 29 380 129 418
rect 29 346 45 380
rect 113 346 129 380
rect 29 330 129 346
rect 187 380 287 418
rect 187 346 203 380
rect 271 346 287 380
rect 187 330 287 346
rect 345 380 445 418
rect 345 346 361 380
rect 429 346 445 380
rect 345 330 445 346
rect 503 380 603 418
rect 503 346 519 380
rect 587 346 603 380
rect 503 330 603 346
rect 661 380 761 418
rect 661 346 677 380
rect 745 346 761 380
rect 661 330 761 346
rect 819 380 919 418
rect 819 346 835 380
rect 903 346 919 380
rect 819 330 919 346
rect 977 380 1077 418
rect 977 346 993 380
rect 1061 346 1077 380
rect 977 330 1077 346
rect 1135 380 1235 418
rect 1135 346 1151 380
rect 1219 346 1235 380
rect 1135 330 1235 346
rect -1235 272 -1135 288
rect -1235 238 -1219 272
rect -1151 238 -1135 272
rect -1235 200 -1135 238
rect -1077 272 -977 288
rect -1077 238 -1061 272
rect -993 238 -977 272
rect -1077 200 -977 238
rect -919 272 -819 288
rect -919 238 -903 272
rect -835 238 -819 272
rect -919 200 -819 238
rect -761 272 -661 288
rect -761 238 -745 272
rect -677 238 -661 272
rect -761 200 -661 238
rect -603 272 -503 288
rect -603 238 -587 272
rect -519 238 -503 272
rect -603 200 -503 238
rect -445 272 -345 288
rect -445 238 -429 272
rect -361 238 -345 272
rect -445 200 -345 238
rect -287 272 -187 288
rect -287 238 -271 272
rect -203 238 -187 272
rect -287 200 -187 238
rect -129 272 -29 288
rect -129 238 -113 272
rect -45 238 -29 272
rect -129 200 -29 238
rect 29 272 129 288
rect 29 238 45 272
rect 113 238 129 272
rect 29 200 129 238
rect 187 272 287 288
rect 187 238 203 272
rect 271 238 287 272
rect 187 200 287 238
rect 345 272 445 288
rect 345 238 361 272
rect 429 238 445 272
rect 345 200 445 238
rect 503 272 603 288
rect 503 238 519 272
rect 587 238 603 272
rect 503 200 603 238
rect 661 272 761 288
rect 661 238 677 272
rect 745 238 761 272
rect 661 200 761 238
rect 819 272 919 288
rect 819 238 835 272
rect 903 238 919 272
rect 819 200 919 238
rect 977 272 1077 288
rect 977 238 993 272
rect 1061 238 1077 272
rect 977 200 1077 238
rect 1135 272 1235 288
rect 1135 238 1151 272
rect 1219 238 1235 272
rect 1135 200 1235 238
rect -1235 -238 -1135 -200
rect -1235 -272 -1219 -238
rect -1151 -272 -1135 -238
rect -1235 -288 -1135 -272
rect -1077 -238 -977 -200
rect -1077 -272 -1061 -238
rect -993 -272 -977 -238
rect -1077 -288 -977 -272
rect -919 -238 -819 -200
rect -919 -272 -903 -238
rect -835 -272 -819 -238
rect -919 -288 -819 -272
rect -761 -238 -661 -200
rect -761 -272 -745 -238
rect -677 -272 -661 -238
rect -761 -288 -661 -272
rect -603 -238 -503 -200
rect -603 -272 -587 -238
rect -519 -272 -503 -238
rect -603 -288 -503 -272
rect -445 -238 -345 -200
rect -445 -272 -429 -238
rect -361 -272 -345 -238
rect -445 -288 -345 -272
rect -287 -238 -187 -200
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -287 -288 -187 -272
rect -129 -238 -29 -200
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect -129 -288 -29 -272
rect 29 -238 129 -200
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 29 -288 129 -272
rect 187 -238 287 -200
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 187 -288 287 -272
rect 345 -238 445 -200
rect 345 -272 361 -238
rect 429 -272 445 -238
rect 345 -288 445 -272
rect 503 -238 603 -200
rect 503 -272 519 -238
rect 587 -272 603 -238
rect 503 -288 603 -272
rect 661 -238 761 -200
rect 661 -272 677 -238
rect 745 -272 761 -238
rect 661 -288 761 -272
rect 819 -238 919 -200
rect 819 -272 835 -238
rect 903 -272 919 -238
rect 819 -288 919 -272
rect 977 -238 1077 -200
rect 977 -272 993 -238
rect 1061 -272 1077 -238
rect 977 -288 1077 -272
rect 1135 -238 1235 -200
rect 1135 -272 1151 -238
rect 1219 -272 1235 -238
rect 1135 -288 1235 -272
rect -1235 -346 -1135 -330
rect -1235 -380 -1219 -346
rect -1151 -380 -1135 -346
rect -1235 -418 -1135 -380
rect -1077 -346 -977 -330
rect -1077 -380 -1061 -346
rect -993 -380 -977 -346
rect -1077 -418 -977 -380
rect -919 -346 -819 -330
rect -919 -380 -903 -346
rect -835 -380 -819 -346
rect -919 -418 -819 -380
rect -761 -346 -661 -330
rect -761 -380 -745 -346
rect -677 -380 -661 -346
rect -761 -418 -661 -380
rect -603 -346 -503 -330
rect -603 -380 -587 -346
rect -519 -380 -503 -346
rect -603 -418 -503 -380
rect -445 -346 -345 -330
rect -445 -380 -429 -346
rect -361 -380 -345 -346
rect -445 -418 -345 -380
rect -287 -346 -187 -330
rect -287 -380 -271 -346
rect -203 -380 -187 -346
rect -287 -418 -187 -380
rect -129 -346 -29 -330
rect -129 -380 -113 -346
rect -45 -380 -29 -346
rect -129 -418 -29 -380
rect 29 -346 129 -330
rect 29 -380 45 -346
rect 113 -380 129 -346
rect 29 -418 129 -380
rect 187 -346 287 -330
rect 187 -380 203 -346
rect 271 -380 287 -346
rect 187 -418 287 -380
rect 345 -346 445 -330
rect 345 -380 361 -346
rect 429 -380 445 -346
rect 345 -418 445 -380
rect 503 -346 603 -330
rect 503 -380 519 -346
rect 587 -380 603 -346
rect 503 -418 603 -380
rect 661 -346 761 -330
rect 661 -380 677 -346
rect 745 -380 761 -346
rect 661 -418 761 -380
rect 819 -346 919 -330
rect 819 -380 835 -346
rect 903 -380 919 -346
rect 819 -418 919 -380
rect 977 -346 1077 -330
rect 977 -380 993 -346
rect 1061 -380 1077 -346
rect 977 -418 1077 -380
rect 1135 -346 1235 -330
rect 1135 -380 1151 -346
rect 1219 -380 1235 -346
rect 1135 -418 1235 -380
rect -1235 -856 -1135 -818
rect -1235 -890 -1219 -856
rect -1151 -890 -1135 -856
rect -1235 -906 -1135 -890
rect -1077 -856 -977 -818
rect -1077 -890 -1061 -856
rect -993 -890 -977 -856
rect -1077 -906 -977 -890
rect -919 -856 -819 -818
rect -919 -890 -903 -856
rect -835 -890 -819 -856
rect -919 -906 -819 -890
rect -761 -856 -661 -818
rect -761 -890 -745 -856
rect -677 -890 -661 -856
rect -761 -906 -661 -890
rect -603 -856 -503 -818
rect -603 -890 -587 -856
rect -519 -890 -503 -856
rect -603 -906 -503 -890
rect -445 -856 -345 -818
rect -445 -890 -429 -856
rect -361 -890 -345 -856
rect -445 -906 -345 -890
rect -287 -856 -187 -818
rect -287 -890 -271 -856
rect -203 -890 -187 -856
rect -287 -906 -187 -890
rect -129 -856 -29 -818
rect -129 -890 -113 -856
rect -45 -890 -29 -856
rect -129 -906 -29 -890
rect 29 -856 129 -818
rect 29 -890 45 -856
rect 113 -890 129 -856
rect 29 -906 129 -890
rect 187 -856 287 -818
rect 187 -890 203 -856
rect 271 -890 287 -856
rect 187 -906 287 -890
rect 345 -856 445 -818
rect 345 -890 361 -856
rect 429 -890 445 -856
rect 345 -906 445 -890
rect 503 -856 603 -818
rect 503 -890 519 -856
rect 587 -890 603 -856
rect 503 -906 603 -890
rect 661 -856 761 -818
rect 661 -890 677 -856
rect 745 -890 761 -856
rect 661 -906 761 -890
rect 819 -856 919 -818
rect 819 -890 835 -856
rect 903 -890 919 -856
rect 819 -906 919 -890
rect 977 -856 1077 -818
rect 977 -890 993 -856
rect 1061 -890 1077 -856
rect 977 -906 1077 -890
rect 1135 -856 1235 -818
rect 1135 -890 1151 -856
rect 1219 -890 1235 -856
rect 1135 -906 1235 -890
<< polycont >>
rect -1219 856 -1151 890
rect -1061 856 -993 890
rect -903 856 -835 890
rect -745 856 -677 890
rect -587 856 -519 890
rect -429 856 -361 890
rect -271 856 -203 890
rect -113 856 -45 890
rect 45 856 113 890
rect 203 856 271 890
rect 361 856 429 890
rect 519 856 587 890
rect 677 856 745 890
rect 835 856 903 890
rect 993 856 1061 890
rect 1151 856 1219 890
rect -1219 346 -1151 380
rect -1061 346 -993 380
rect -903 346 -835 380
rect -745 346 -677 380
rect -587 346 -519 380
rect -429 346 -361 380
rect -271 346 -203 380
rect -113 346 -45 380
rect 45 346 113 380
rect 203 346 271 380
rect 361 346 429 380
rect 519 346 587 380
rect 677 346 745 380
rect 835 346 903 380
rect 993 346 1061 380
rect 1151 346 1219 380
rect -1219 238 -1151 272
rect -1061 238 -993 272
rect -903 238 -835 272
rect -745 238 -677 272
rect -587 238 -519 272
rect -429 238 -361 272
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect 361 238 429 272
rect 519 238 587 272
rect 677 238 745 272
rect 835 238 903 272
rect 993 238 1061 272
rect 1151 238 1219 272
rect -1219 -272 -1151 -238
rect -1061 -272 -993 -238
rect -903 -272 -835 -238
rect -745 -272 -677 -238
rect -587 -272 -519 -238
rect -429 -272 -361 -238
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
rect 361 -272 429 -238
rect 519 -272 587 -238
rect 677 -272 745 -238
rect 835 -272 903 -238
rect 993 -272 1061 -238
rect 1151 -272 1219 -238
rect -1219 -380 -1151 -346
rect -1061 -380 -993 -346
rect -903 -380 -835 -346
rect -745 -380 -677 -346
rect -587 -380 -519 -346
rect -429 -380 -361 -346
rect -271 -380 -203 -346
rect -113 -380 -45 -346
rect 45 -380 113 -346
rect 203 -380 271 -346
rect 361 -380 429 -346
rect 519 -380 587 -346
rect 677 -380 745 -346
rect 835 -380 903 -346
rect 993 -380 1061 -346
rect 1151 -380 1219 -346
rect -1219 -890 -1151 -856
rect -1061 -890 -993 -856
rect -903 -890 -835 -856
rect -745 -890 -677 -856
rect -587 -890 -519 -856
rect -429 -890 -361 -856
rect -271 -890 -203 -856
rect -113 -890 -45 -856
rect 45 -890 113 -856
rect 203 -890 271 -856
rect 361 -890 429 -856
rect 519 -890 587 -856
rect 677 -890 745 -856
rect 835 -890 903 -856
rect 993 -890 1061 -856
rect 1151 -890 1219 -856
<< locali >>
rect -1395 958 -1299 992
rect 1299 958 1395 992
rect -1395 896 -1361 958
rect 1361 896 1395 958
rect -1235 856 -1219 890
rect -1151 856 -1135 890
rect -1077 856 -1061 890
rect -993 856 -977 890
rect -919 856 -903 890
rect -835 856 -819 890
rect -761 856 -745 890
rect -677 856 -661 890
rect -603 856 -587 890
rect -519 856 -503 890
rect -445 856 -429 890
rect -361 856 -345 890
rect -287 856 -271 890
rect -203 856 -187 890
rect -129 856 -113 890
rect -45 856 -29 890
rect 29 856 45 890
rect 113 856 129 890
rect 187 856 203 890
rect 271 856 287 890
rect 345 856 361 890
rect 429 856 445 890
rect 503 856 519 890
rect 587 856 603 890
rect 661 856 677 890
rect 745 856 761 890
rect 819 856 835 890
rect 903 856 919 890
rect 977 856 993 890
rect 1061 856 1077 890
rect 1135 856 1151 890
rect 1219 856 1235 890
rect -1281 806 -1247 822
rect -1281 414 -1247 430
rect -1123 806 -1089 822
rect -1123 414 -1089 430
rect -965 806 -931 822
rect -965 414 -931 430
rect -807 806 -773 822
rect -807 414 -773 430
rect -649 806 -615 822
rect -649 414 -615 430
rect -491 806 -457 822
rect -491 414 -457 430
rect -333 806 -299 822
rect -333 414 -299 430
rect -175 806 -141 822
rect -175 414 -141 430
rect -17 806 17 822
rect -17 414 17 430
rect 141 806 175 822
rect 141 414 175 430
rect 299 806 333 822
rect 299 414 333 430
rect 457 806 491 822
rect 457 414 491 430
rect 615 806 649 822
rect 615 414 649 430
rect 773 806 807 822
rect 773 414 807 430
rect 931 806 965 822
rect 931 414 965 430
rect 1089 806 1123 822
rect 1089 414 1123 430
rect 1247 806 1281 822
rect 1247 414 1281 430
rect -1235 346 -1219 380
rect -1151 346 -1135 380
rect -1077 346 -1061 380
rect -993 346 -977 380
rect -919 346 -903 380
rect -835 346 -819 380
rect -761 346 -745 380
rect -677 346 -661 380
rect -603 346 -587 380
rect -519 346 -503 380
rect -445 346 -429 380
rect -361 346 -345 380
rect -287 346 -271 380
rect -203 346 -187 380
rect -129 346 -113 380
rect -45 346 -29 380
rect 29 346 45 380
rect 113 346 129 380
rect 187 346 203 380
rect 271 346 287 380
rect 345 346 361 380
rect 429 346 445 380
rect 503 346 519 380
rect 587 346 603 380
rect 661 346 677 380
rect 745 346 761 380
rect 819 346 835 380
rect 903 346 919 380
rect 977 346 993 380
rect 1061 346 1077 380
rect 1135 346 1151 380
rect 1219 346 1235 380
rect -1235 238 -1219 272
rect -1151 238 -1135 272
rect -1077 238 -1061 272
rect -993 238 -977 272
rect -919 238 -903 272
rect -835 238 -819 272
rect -761 238 -745 272
rect -677 238 -661 272
rect -603 238 -587 272
rect -519 238 -503 272
rect -445 238 -429 272
rect -361 238 -345 272
rect -287 238 -271 272
rect -203 238 -187 272
rect -129 238 -113 272
rect -45 238 -29 272
rect 29 238 45 272
rect 113 238 129 272
rect 187 238 203 272
rect 271 238 287 272
rect 345 238 361 272
rect 429 238 445 272
rect 503 238 519 272
rect 587 238 603 272
rect 661 238 677 272
rect 745 238 761 272
rect 819 238 835 272
rect 903 238 919 272
rect 977 238 993 272
rect 1061 238 1077 272
rect 1135 238 1151 272
rect 1219 238 1235 272
rect -1281 188 -1247 204
rect -1281 -204 -1247 -188
rect -1123 188 -1089 204
rect -1123 -204 -1089 -188
rect -965 188 -931 204
rect -965 -204 -931 -188
rect -807 188 -773 204
rect -807 -204 -773 -188
rect -649 188 -615 204
rect -649 -204 -615 -188
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect 615 188 649 204
rect 615 -204 649 -188
rect 773 188 807 204
rect 773 -204 807 -188
rect 931 188 965 204
rect 931 -204 965 -188
rect 1089 188 1123 204
rect 1089 -204 1123 -188
rect 1247 188 1281 204
rect 1247 -204 1281 -188
rect -1235 -272 -1219 -238
rect -1151 -272 -1135 -238
rect -1077 -272 -1061 -238
rect -993 -272 -977 -238
rect -919 -272 -903 -238
rect -835 -272 -819 -238
rect -761 -272 -745 -238
rect -677 -272 -661 -238
rect -603 -272 -587 -238
rect -519 -272 -503 -238
rect -445 -272 -429 -238
rect -361 -272 -345 -238
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 345 -272 361 -238
rect 429 -272 445 -238
rect 503 -272 519 -238
rect 587 -272 603 -238
rect 661 -272 677 -238
rect 745 -272 761 -238
rect 819 -272 835 -238
rect 903 -272 919 -238
rect 977 -272 993 -238
rect 1061 -272 1077 -238
rect 1135 -272 1151 -238
rect 1219 -272 1235 -238
rect -1235 -380 -1219 -346
rect -1151 -380 -1135 -346
rect -1077 -380 -1061 -346
rect -993 -380 -977 -346
rect -919 -380 -903 -346
rect -835 -380 -819 -346
rect -761 -380 -745 -346
rect -677 -380 -661 -346
rect -603 -380 -587 -346
rect -519 -380 -503 -346
rect -445 -380 -429 -346
rect -361 -380 -345 -346
rect -287 -380 -271 -346
rect -203 -380 -187 -346
rect -129 -380 -113 -346
rect -45 -380 -29 -346
rect 29 -380 45 -346
rect 113 -380 129 -346
rect 187 -380 203 -346
rect 271 -380 287 -346
rect 345 -380 361 -346
rect 429 -380 445 -346
rect 503 -380 519 -346
rect 587 -380 603 -346
rect 661 -380 677 -346
rect 745 -380 761 -346
rect 819 -380 835 -346
rect 903 -380 919 -346
rect 977 -380 993 -346
rect 1061 -380 1077 -346
rect 1135 -380 1151 -346
rect 1219 -380 1235 -346
rect -1281 -430 -1247 -414
rect -1281 -822 -1247 -806
rect -1123 -430 -1089 -414
rect -1123 -822 -1089 -806
rect -965 -430 -931 -414
rect -965 -822 -931 -806
rect -807 -430 -773 -414
rect -807 -822 -773 -806
rect -649 -430 -615 -414
rect -649 -822 -615 -806
rect -491 -430 -457 -414
rect -491 -822 -457 -806
rect -333 -430 -299 -414
rect -333 -822 -299 -806
rect -175 -430 -141 -414
rect -175 -822 -141 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 141 -430 175 -414
rect 141 -822 175 -806
rect 299 -430 333 -414
rect 299 -822 333 -806
rect 457 -430 491 -414
rect 457 -822 491 -806
rect 615 -430 649 -414
rect 615 -822 649 -806
rect 773 -430 807 -414
rect 773 -822 807 -806
rect 931 -430 965 -414
rect 931 -822 965 -806
rect 1089 -430 1123 -414
rect 1089 -822 1123 -806
rect 1247 -430 1281 -414
rect 1247 -822 1281 -806
rect -1235 -890 -1219 -856
rect -1151 -890 -1135 -856
rect -1077 -890 -1061 -856
rect -993 -890 -977 -856
rect -919 -890 -903 -856
rect -835 -890 -819 -856
rect -761 -890 -745 -856
rect -677 -890 -661 -856
rect -603 -890 -587 -856
rect -519 -890 -503 -856
rect -445 -890 -429 -856
rect -361 -890 -345 -856
rect -287 -890 -271 -856
rect -203 -890 -187 -856
rect -129 -890 -113 -856
rect -45 -890 -29 -856
rect 29 -890 45 -856
rect 113 -890 129 -856
rect 187 -890 203 -856
rect 271 -890 287 -856
rect 345 -890 361 -856
rect 429 -890 445 -856
rect 503 -890 519 -856
rect 587 -890 603 -856
rect 661 -890 677 -856
rect 745 -890 761 -856
rect 819 -890 835 -856
rect 903 -890 919 -856
rect 977 -890 993 -856
rect 1061 -890 1077 -856
rect 1135 -890 1151 -856
rect 1219 -890 1235 -856
rect -1395 -958 -1361 -896
rect 1361 -958 1395 -896
rect -1395 -992 -1299 -958
rect 1299 -992 1395 -958
<< viali >>
rect -1219 856 -1151 890
rect -1061 856 -993 890
rect -903 856 -835 890
rect -745 856 -677 890
rect -587 856 -519 890
rect -429 856 -361 890
rect -271 856 -203 890
rect -113 856 -45 890
rect 45 856 113 890
rect 203 856 271 890
rect 361 856 429 890
rect 519 856 587 890
rect 677 856 745 890
rect 835 856 903 890
rect 993 856 1061 890
rect 1151 856 1219 890
rect -1281 430 -1247 806
rect -1123 430 -1089 806
rect -965 430 -931 806
rect -807 430 -773 806
rect -649 430 -615 806
rect -491 430 -457 806
rect -333 430 -299 806
rect -175 430 -141 806
rect -17 430 17 806
rect 141 430 175 806
rect 299 430 333 806
rect 457 430 491 806
rect 615 430 649 806
rect 773 430 807 806
rect 931 430 965 806
rect 1089 430 1123 806
rect 1247 430 1281 806
rect -1219 346 -1151 380
rect -1061 346 -993 380
rect -903 346 -835 380
rect -745 346 -677 380
rect -587 346 -519 380
rect -429 346 -361 380
rect -271 346 -203 380
rect -113 346 -45 380
rect 45 346 113 380
rect 203 346 271 380
rect 361 346 429 380
rect 519 346 587 380
rect 677 346 745 380
rect 835 346 903 380
rect 993 346 1061 380
rect 1151 346 1219 380
rect -1219 238 -1151 272
rect -1061 238 -993 272
rect -903 238 -835 272
rect -745 238 -677 272
rect -587 238 -519 272
rect -429 238 -361 272
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect 361 238 429 272
rect 519 238 587 272
rect 677 238 745 272
rect 835 238 903 272
rect 993 238 1061 272
rect 1151 238 1219 272
rect -1281 -188 -1247 188
rect -1123 -188 -1089 188
rect -965 -188 -931 188
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect 931 -188 965 188
rect 1089 -188 1123 188
rect 1247 -188 1281 188
rect -1219 -272 -1151 -238
rect -1061 -272 -993 -238
rect -903 -272 -835 -238
rect -745 -272 -677 -238
rect -587 -272 -519 -238
rect -429 -272 -361 -238
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
rect 361 -272 429 -238
rect 519 -272 587 -238
rect 677 -272 745 -238
rect 835 -272 903 -238
rect 993 -272 1061 -238
rect 1151 -272 1219 -238
rect -1219 -380 -1151 -346
rect -1061 -380 -993 -346
rect -903 -380 -835 -346
rect -745 -380 -677 -346
rect -587 -380 -519 -346
rect -429 -380 -361 -346
rect -271 -380 -203 -346
rect -113 -380 -45 -346
rect 45 -380 113 -346
rect 203 -380 271 -346
rect 361 -380 429 -346
rect 519 -380 587 -346
rect 677 -380 745 -346
rect 835 -380 903 -346
rect 993 -380 1061 -346
rect 1151 -380 1219 -346
rect -1281 -806 -1247 -430
rect -1123 -806 -1089 -430
rect -965 -806 -931 -430
rect -807 -806 -773 -430
rect -649 -806 -615 -430
rect -491 -806 -457 -430
rect -333 -806 -299 -430
rect -175 -806 -141 -430
rect -17 -806 17 -430
rect 141 -806 175 -430
rect 299 -806 333 -430
rect 457 -806 491 -430
rect 615 -806 649 -430
rect 773 -806 807 -430
rect 931 -806 965 -430
rect 1089 -806 1123 -430
rect 1247 -806 1281 -430
rect -1219 -890 -1151 -856
rect -1061 -890 -993 -856
rect -903 -890 -835 -856
rect -745 -890 -677 -856
rect -587 -890 -519 -856
rect -429 -890 -361 -856
rect -271 -890 -203 -856
rect -113 -890 -45 -856
rect 45 -890 113 -856
rect 203 -890 271 -856
rect 361 -890 429 -856
rect 519 -890 587 -856
rect 677 -890 745 -856
rect 835 -890 903 -856
rect 993 -890 1061 -856
rect 1151 -890 1219 -856
<< metal1 >>
rect -1231 890 -1139 896
rect -1231 856 -1219 890
rect -1151 856 -1139 890
rect -1231 850 -1139 856
rect -1073 890 -981 896
rect -1073 856 -1061 890
rect -993 856 -981 890
rect -1073 850 -981 856
rect -915 890 -823 896
rect -915 856 -903 890
rect -835 856 -823 890
rect -915 850 -823 856
rect -757 890 -665 896
rect -757 856 -745 890
rect -677 856 -665 890
rect -757 850 -665 856
rect -599 890 -507 896
rect -599 856 -587 890
rect -519 856 -507 890
rect -599 850 -507 856
rect -441 890 -349 896
rect -441 856 -429 890
rect -361 856 -349 890
rect -441 850 -349 856
rect -283 890 -191 896
rect -283 856 -271 890
rect -203 856 -191 890
rect -283 850 -191 856
rect -125 890 -33 896
rect -125 856 -113 890
rect -45 856 -33 890
rect -125 850 -33 856
rect 33 890 125 896
rect 33 856 45 890
rect 113 856 125 890
rect 33 850 125 856
rect 191 890 283 896
rect 191 856 203 890
rect 271 856 283 890
rect 191 850 283 856
rect 349 890 441 896
rect 349 856 361 890
rect 429 856 441 890
rect 349 850 441 856
rect 507 890 599 896
rect 507 856 519 890
rect 587 856 599 890
rect 507 850 599 856
rect 665 890 757 896
rect 665 856 677 890
rect 745 856 757 890
rect 665 850 757 856
rect 823 890 915 896
rect 823 856 835 890
rect 903 856 915 890
rect 823 850 915 856
rect 981 890 1073 896
rect 981 856 993 890
rect 1061 856 1073 890
rect 981 850 1073 856
rect 1139 890 1231 896
rect 1139 856 1151 890
rect 1219 856 1231 890
rect 1139 850 1231 856
rect -1287 806 -1241 818
rect -1287 430 -1281 806
rect -1247 430 -1241 806
rect -1287 418 -1241 430
rect -1129 806 -1083 818
rect -1129 430 -1123 806
rect -1089 430 -1083 806
rect -1129 418 -1083 430
rect -971 806 -925 818
rect -971 430 -965 806
rect -931 430 -925 806
rect -971 418 -925 430
rect -813 806 -767 818
rect -813 430 -807 806
rect -773 430 -767 806
rect -813 418 -767 430
rect -655 806 -609 818
rect -655 430 -649 806
rect -615 430 -609 806
rect -655 418 -609 430
rect -497 806 -451 818
rect -497 430 -491 806
rect -457 430 -451 806
rect -497 418 -451 430
rect -339 806 -293 818
rect -339 430 -333 806
rect -299 430 -293 806
rect -339 418 -293 430
rect -181 806 -135 818
rect -181 430 -175 806
rect -141 430 -135 806
rect -181 418 -135 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 135 806 181 818
rect 135 430 141 806
rect 175 430 181 806
rect 135 418 181 430
rect 293 806 339 818
rect 293 430 299 806
rect 333 430 339 806
rect 293 418 339 430
rect 451 806 497 818
rect 451 430 457 806
rect 491 430 497 806
rect 451 418 497 430
rect 609 806 655 818
rect 609 430 615 806
rect 649 430 655 806
rect 609 418 655 430
rect 767 806 813 818
rect 767 430 773 806
rect 807 430 813 806
rect 767 418 813 430
rect 925 806 971 818
rect 925 430 931 806
rect 965 430 971 806
rect 925 418 971 430
rect 1083 806 1129 818
rect 1083 430 1089 806
rect 1123 430 1129 806
rect 1083 418 1129 430
rect 1241 806 1287 818
rect 1241 430 1247 806
rect 1281 430 1287 806
rect 1241 418 1287 430
rect -1231 380 -1139 386
rect -1231 346 -1219 380
rect -1151 346 -1139 380
rect -1231 340 -1139 346
rect -1073 380 -981 386
rect -1073 346 -1061 380
rect -993 346 -981 380
rect -1073 340 -981 346
rect -915 380 -823 386
rect -915 346 -903 380
rect -835 346 -823 380
rect -915 340 -823 346
rect -757 380 -665 386
rect -757 346 -745 380
rect -677 346 -665 380
rect -757 340 -665 346
rect -599 380 -507 386
rect -599 346 -587 380
rect -519 346 -507 380
rect -599 340 -507 346
rect -441 380 -349 386
rect -441 346 -429 380
rect -361 346 -349 380
rect -441 340 -349 346
rect -283 380 -191 386
rect -283 346 -271 380
rect -203 346 -191 380
rect -283 340 -191 346
rect -125 380 -33 386
rect -125 346 -113 380
rect -45 346 -33 380
rect -125 340 -33 346
rect 33 380 125 386
rect 33 346 45 380
rect 113 346 125 380
rect 33 340 125 346
rect 191 380 283 386
rect 191 346 203 380
rect 271 346 283 380
rect 191 340 283 346
rect 349 380 441 386
rect 349 346 361 380
rect 429 346 441 380
rect 349 340 441 346
rect 507 380 599 386
rect 507 346 519 380
rect 587 346 599 380
rect 507 340 599 346
rect 665 380 757 386
rect 665 346 677 380
rect 745 346 757 380
rect 665 340 757 346
rect 823 380 915 386
rect 823 346 835 380
rect 903 346 915 380
rect 823 340 915 346
rect 981 380 1073 386
rect 981 346 993 380
rect 1061 346 1073 380
rect 981 340 1073 346
rect 1139 380 1231 386
rect 1139 346 1151 380
rect 1219 346 1231 380
rect 1139 340 1231 346
rect -1231 272 -1139 278
rect -1231 238 -1219 272
rect -1151 238 -1139 272
rect -1231 232 -1139 238
rect -1073 272 -981 278
rect -1073 238 -1061 272
rect -993 238 -981 272
rect -1073 232 -981 238
rect -915 272 -823 278
rect -915 238 -903 272
rect -835 238 -823 272
rect -915 232 -823 238
rect -757 272 -665 278
rect -757 238 -745 272
rect -677 238 -665 272
rect -757 232 -665 238
rect -599 272 -507 278
rect -599 238 -587 272
rect -519 238 -507 272
rect -599 232 -507 238
rect -441 272 -349 278
rect -441 238 -429 272
rect -361 238 -349 272
rect -441 232 -349 238
rect -283 272 -191 278
rect -283 238 -271 272
rect -203 238 -191 272
rect -283 232 -191 238
rect -125 272 -33 278
rect -125 238 -113 272
rect -45 238 -33 272
rect -125 232 -33 238
rect 33 272 125 278
rect 33 238 45 272
rect 113 238 125 272
rect 33 232 125 238
rect 191 272 283 278
rect 191 238 203 272
rect 271 238 283 272
rect 191 232 283 238
rect 349 272 441 278
rect 349 238 361 272
rect 429 238 441 272
rect 349 232 441 238
rect 507 272 599 278
rect 507 238 519 272
rect 587 238 599 272
rect 507 232 599 238
rect 665 272 757 278
rect 665 238 677 272
rect 745 238 757 272
rect 665 232 757 238
rect 823 272 915 278
rect 823 238 835 272
rect 903 238 915 272
rect 823 232 915 238
rect 981 272 1073 278
rect 981 238 993 272
rect 1061 238 1073 272
rect 981 232 1073 238
rect 1139 272 1231 278
rect 1139 238 1151 272
rect 1219 238 1231 272
rect 1139 232 1231 238
rect -1287 188 -1241 200
rect -1287 -188 -1281 188
rect -1247 -188 -1241 188
rect -1287 -200 -1241 -188
rect -1129 188 -1083 200
rect -1129 -188 -1123 188
rect -1089 -188 -1083 188
rect -1129 -200 -1083 -188
rect -971 188 -925 200
rect -971 -188 -965 188
rect -931 -188 -925 188
rect -971 -200 -925 -188
rect -813 188 -767 200
rect -813 -188 -807 188
rect -773 -188 -767 188
rect -813 -200 -767 -188
rect -655 188 -609 200
rect -655 -188 -649 188
rect -615 -188 -609 188
rect -655 -200 -609 -188
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect 609 188 655 200
rect 609 -188 615 188
rect 649 -188 655 188
rect 609 -200 655 -188
rect 767 188 813 200
rect 767 -188 773 188
rect 807 -188 813 188
rect 767 -200 813 -188
rect 925 188 971 200
rect 925 -188 931 188
rect 965 -188 971 188
rect 925 -200 971 -188
rect 1083 188 1129 200
rect 1083 -188 1089 188
rect 1123 -188 1129 188
rect 1083 -200 1129 -188
rect 1241 188 1287 200
rect 1241 -188 1247 188
rect 1281 -188 1287 188
rect 1241 -200 1287 -188
rect -1231 -238 -1139 -232
rect -1231 -272 -1219 -238
rect -1151 -272 -1139 -238
rect -1231 -278 -1139 -272
rect -1073 -238 -981 -232
rect -1073 -272 -1061 -238
rect -993 -272 -981 -238
rect -1073 -278 -981 -272
rect -915 -238 -823 -232
rect -915 -272 -903 -238
rect -835 -272 -823 -238
rect -915 -278 -823 -272
rect -757 -238 -665 -232
rect -757 -272 -745 -238
rect -677 -272 -665 -238
rect -757 -278 -665 -272
rect -599 -238 -507 -232
rect -599 -272 -587 -238
rect -519 -272 -507 -238
rect -599 -278 -507 -272
rect -441 -238 -349 -232
rect -441 -272 -429 -238
rect -361 -272 -349 -238
rect -441 -278 -349 -272
rect -283 -238 -191 -232
rect -283 -272 -271 -238
rect -203 -272 -191 -238
rect -283 -278 -191 -272
rect -125 -238 -33 -232
rect -125 -272 -113 -238
rect -45 -272 -33 -238
rect -125 -278 -33 -272
rect 33 -238 125 -232
rect 33 -272 45 -238
rect 113 -272 125 -238
rect 33 -278 125 -272
rect 191 -238 283 -232
rect 191 -272 203 -238
rect 271 -272 283 -238
rect 191 -278 283 -272
rect 349 -238 441 -232
rect 349 -272 361 -238
rect 429 -272 441 -238
rect 349 -278 441 -272
rect 507 -238 599 -232
rect 507 -272 519 -238
rect 587 -272 599 -238
rect 507 -278 599 -272
rect 665 -238 757 -232
rect 665 -272 677 -238
rect 745 -272 757 -238
rect 665 -278 757 -272
rect 823 -238 915 -232
rect 823 -272 835 -238
rect 903 -272 915 -238
rect 823 -278 915 -272
rect 981 -238 1073 -232
rect 981 -272 993 -238
rect 1061 -272 1073 -238
rect 981 -278 1073 -272
rect 1139 -238 1231 -232
rect 1139 -272 1151 -238
rect 1219 -272 1231 -238
rect 1139 -278 1231 -272
rect -1231 -346 -1139 -340
rect -1231 -380 -1219 -346
rect -1151 -380 -1139 -346
rect -1231 -386 -1139 -380
rect -1073 -346 -981 -340
rect -1073 -380 -1061 -346
rect -993 -380 -981 -346
rect -1073 -386 -981 -380
rect -915 -346 -823 -340
rect -915 -380 -903 -346
rect -835 -380 -823 -346
rect -915 -386 -823 -380
rect -757 -346 -665 -340
rect -757 -380 -745 -346
rect -677 -380 -665 -346
rect -757 -386 -665 -380
rect -599 -346 -507 -340
rect -599 -380 -587 -346
rect -519 -380 -507 -346
rect -599 -386 -507 -380
rect -441 -346 -349 -340
rect -441 -380 -429 -346
rect -361 -380 -349 -346
rect -441 -386 -349 -380
rect -283 -346 -191 -340
rect -283 -380 -271 -346
rect -203 -380 -191 -346
rect -283 -386 -191 -380
rect -125 -346 -33 -340
rect -125 -380 -113 -346
rect -45 -380 -33 -346
rect -125 -386 -33 -380
rect 33 -346 125 -340
rect 33 -380 45 -346
rect 113 -380 125 -346
rect 33 -386 125 -380
rect 191 -346 283 -340
rect 191 -380 203 -346
rect 271 -380 283 -346
rect 191 -386 283 -380
rect 349 -346 441 -340
rect 349 -380 361 -346
rect 429 -380 441 -346
rect 349 -386 441 -380
rect 507 -346 599 -340
rect 507 -380 519 -346
rect 587 -380 599 -346
rect 507 -386 599 -380
rect 665 -346 757 -340
rect 665 -380 677 -346
rect 745 -380 757 -346
rect 665 -386 757 -380
rect 823 -346 915 -340
rect 823 -380 835 -346
rect 903 -380 915 -346
rect 823 -386 915 -380
rect 981 -346 1073 -340
rect 981 -380 993 -346
rect 1061 -380 1073 -346
rect 981 -386 1073 -380
rect 1139 -346 1231 -340
rect 1139 -380 1151 -346
rect 1219 -380 1231 -346
rect 1139 -386 1231 -380
rect -1287 -430 -1241 -418
rect -1287 -806 -1281 -430
rect -1247 -806 -1241 -430
rect -1287 -818 -1241 -806
rect -1129 -430 -1083 -418
rect -1129 -806 -1123 -430
rect -1089 -806 -1083 -430
rect -1129 -818 -1083 -806
rect -971 -430 -925 -418
rect -971 -806 -965 -430
rect -931 -806 -925 -430
rect -971 -818 -925 -806
rect -813 -430 -767 -418
rect -813 -806 -807 -430
rect -773 -806 -767 -430
rect -813 -818 -767 -806
rect -655 -430 -609 -418
rect -655 -806 -649 -430
rect -615 -806 -609 -430
rect -655 -818 -609 -806
rect -497 -430 -451 -418
rect -497 -806 -491 -430
rect -457 -806 -451 -430
rect -497 -818 -451 -806
rect -339 -430 -293 -418
rect -339 -806 -333 -430
rect -299 -806 -293 -430
rect -339 -818 -293 -806
rect -181 -430 -135 -418
rect -181 -806 -175 -430
rect -141 -806 -135 -430
rect -181 -818 -135 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 135 -430 181 -418
rect 135 -806 141 -430
rect 175 -806 181 -430
rect 135 -818 181 -806
rect 293 -430 339 -418
rect 293 -806 299 -430
rect 333 -806 339 -430
rect 293 -818 339 -806
rect 451 -430 497 -418
rect 451 -806 457 -430
rect 491 -806 497 -430
rect 451 -818 497 -806
rect 609 -430 655 -418
rect 609 -806 615 -430
rect 649 -806 655 -430
rect 609 -818 655 -806
rect 767 -430 813 -418
rect 767 -806 773 -430
rect 807 -806 813 -430
rect 767 -818 813 -806
rect 925 -430 971 -418
rect 925 -806 931 -430
rect 965 -806 971 -430
rect 925 -818 971 -806
rect 1083 -430 1129 -418
rect 1083 -806 1089 -430
rect 1123 -806 1129 -430
rect 1083 -818 1129 -806
rect 1241 -430 1287 -418
rect 1241 -806 1247 -430
rect 1281 -806 1287 -430
rect 1241 -818 1287 -806
rect -1231 -856 -1139 -850
rect -1231 -890 -1219 -856
rect -1151 -890 -1139 -856
rect -1231 -896 -1139 -890
rect -1073 -856 -981 -850
rect -1073 -890 -1061 -856
rect -993 -890 -981 -856
rect -1073 -896 -981 -890
rect -915 -856 -823 -850
rect -915 -890 -903 -856
rect -835 -890 -823 -856
rect -915 -896 -823 -890
rect -757 -856 -665 -850
rect -757 -890 -745 -856
rect -677 -890 -665 -856
rect -757 -896 -665 -890
rect -599 -856 -507 -850
rect -599 -890 -587 -856
rect -519 -890 -507 -856
rect -599 -896 -507 -890
rect -441 -856 -349 -850
rect -441 -890 -429 -856
rect -361 -890 -349 -856
rect -441 -896 -349 -890
rect -283 -856 -191 -850
rect -283 -890 -271 -856
rect -203 -890 -191 -856
rect -283 -896 -191 -890
rect -125 -856 -33 -850
rect -125 -890 -113 -856
rect -45 -890 -33 -856
rect -125 -896 -33 -890
rect 33 -856 125 -850
rect 33 -890 45 -856
rect 113 -890 125 -856
rect 33 -896 125 -890
rect 191 -856 283 -850
rect 191 -890 203 -856
rect 271 -890 283 -856
rect 191 -896 283 -890
rect 349 -856 441 -850
rect 349 -890 361 -856
rect 429 -890 441 -856
rect 349 -896 441 -890
rect 507 -856 599 -850
rect 507 -890 519 -856
rect 587 -890 599 -856
rect 507 -896 599 -890
rect 665 -856 757 -850
rect 665 -890 677 -856
rect 745 -890 757 -856
rect 665 -896 757 -890
rect 823 -856 915 -850
rect 823 -890 835 -856
rect 903 -890 915 -856
rect 823 -896 915 -890
rect 981 -856 1073 -850
rect 981 -890 993 -856
rect 1061 -890 1073 -856
rect 981 -896 1073 -890
rect 1139 -856 1231 -850
rect 1139 -890 1151 -856
rect 1219 -890 1231 -856
rect 1139 -896 1231 -890
<< properties >>
string FIXED_BBOX -1378 -975 1378 975
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.5 m 3 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
