magic
tech sky130B
magscale 1 2
timestamp 1654606386
<< error_p >>
rect -2141 599 -2083 605
rect -1949 599 -1891 605
rect -1757 599 -1699 605
rect -1565 599 -1507 605
rect -1373 599 -1315 605
rect -1181 599 -1123 605
rect -989 599 -931 605
rect -797 599 -739 605
rect -605 599 -547 605
rect -413 599 -355 605
rect -221 599 -163 605
rect -29 599 29 605
rect 163 599 221 605
rect 355 599 413 605
rect 547 599 605 605
rect 739 599 797 605
rect 931 599 989 605
rect 1123 599 1181 605
rect 1315 599 1373 605
rect 1507 599 1565 605
rect 1699 599 1757 605
rect 1891 599 1949 605
rect 2083 599 2141 605
rect -2141 565 -2129 599
rect -1949 565 -1937 599
rect -1757 565 -1745 599
rect -1565 565 -1553 599
rect -1373 565 -1361 599
rect -1181 565 -1169 599
rect -989 565 -977 599
rect -797 565 -785 599
rect -605 565 -593 599
rect -413 565 -401 599
rect -221 565 -209 599
rect -29 565 -17 599
rect 163 565 175 599
rect 355 565 367 599
rect 547 565 559 599
rect 739 565 751 599
rect 931 565 943 599
rect 1123 565 1135 599
rect 1315 565 1327 599
rect 1507 565 1519 599
rect 1699 565 1711 599
rect 1891 565 1903 599
rect 2083 565 2095 599
rect -2141 559 -2083 565
rect -1949 559 -1891 565
rect -1757 559 -1699 565
rect -1565 559 -1507 565
rect -1373 559 -1315 565
rect -1181 559 -1123 565
rect -989 559 -931 565
rect -797 559 -739 565
rect -605 559 -547 565
rect -413 559 -355 565
rect -221 559 -163 565
rect -29 559 29 565
rect 163 559 221 565
rect 355 559 413 565
rect 547 559 605 565
rect 739 559 797 565
rect 931 559 989 565
rect 1123 559 1181 565
rect 1315 559 1373 565
rect 1507 559 1565 565
rect 1699 559 1757 565
rect 1891 559 1949 565
rect 2083 559 2141 565
rect -2045 71 -1987 77
rect -1853 71 -1795 77
rect -1661 71 -1603 77
rect -1469 71 -1411 77
rect -1277 71 -1219 77
rect -1085 71 -1027 77
rect -893 71 -835 77
rect -701 71 -643 77
rect -509 71 -451 77
rect -317 71 -259 77
rect -125 71 -67 77
rect 67 71 125 77
rect 259 71 317 77
rect 451 71 509 77
rect 643 71 701 77
rect 835 71 893 77
rect 1027 71 1085 77
rect 1219 71 1277 77
rect 1411 71 1469 77
rect 1603 71 1661 77
rect 1795 71 1853 77
rect 1987 71 2045 77
rect -2045 37 -2033 71
rect -1853 37 -1841 71
rect -1661 37 -1649 71
rect -1469 37 -1457 71
rect -1277 37 -1265 71
rect -1085 37 -1073 71
rect -893 37 -881 71
rect -701 37 -689 71
rect -509 37 -497 71
rect -317 37 -305 71
rect -125 37 -113 71
rect 67 37 79 71
rect 259 37 271 71
rect 451 37 463 71
rect 643 37 655 71
rect 835 37 847 71
rect 1027 37 1039 71
rect 1219 37 1231 71
rect 1411 37 1423 71
rect 1603 37 1615 71
rect 1795 37 1807 71
rect 1987 37 1999 71
rect -2045 31 -1987 37
rect -1853 31 -1795 37
rect -1661 31 -1603 37
rect -1469 31 -1411 37
rect -1277 31 -1219 37
rect -1085 31 -1027 37
rect -893 31 -835 37
rect -701 31 -643 37
rect -509 31 -451 37
rect -317 31 -259 37
rect -125 31 -67 37
rect 67 31 125 37
rect 259 31 317 37
rect 451 31 509 37
rect 643 31 701 37
rect 835 31 893 37
rect 1027 31 1085 37
rect 1219 31 1277 37
rect 1411 31 1469 37
rect 1603 31 1661 37
rect 1795 31 1853 37
rect 1987 31 2045 37
rect -2045 -37 -1987 -31
rect -1853 -37 -1795 -31
rect -1661 -37 -1603 -31
rect -1469 -37 -1411 -31
rect -1277 -37 -1219 -31
rect -1085 -37 -1027 -31
rect -893 -37 -835 -31
rect -701 -37 -643 -31
rect -509 -37 -451 -31
rect -317 -37 -259 -31
rect -125 -37 -67 -31
rect 67 -37 125 -31
rect 259 -37 317 -31
rect 451 -37 509 -31
rect 643 -37 701 -31
rect 835 -37 893 -31
rect 1027 -37 1085 -31
rect 1219 -37 1277 -31
rect 1411 -37 1469 -31
rect 1603 -37 1661 -31
rect 1795 -37 1853 -31
rect 1987 -37 2045 -31
rect -2045 -71 -2033 -37
rect -1853 -71 -1841 -37
rect -1661 -71 -1649 -37
rect -1469 -71 -1457 -37
rect -1277 -71 -1265 -37
rect -1085 -71 -1073 -37
rect -893 -71 -881 -37
rect -701 -71 -689 -37
rect -509 -71 -497 -37
rect -317 -71 -305 -37
rect -125 -71 -113 -37
rect 67 -71 79 -37
rect 259 -71 271 -37
rect 451 -71 463 -37
rect 643 -71 655 -37
rect 835 -71 847 -37
rect 1027 -71 1039 -37
rect 1219 -71 1231 -37
rect 1411 -71 1423 -37
rect 1603 -71 1615 -37
rect 1795 -71 1807 -37
rect 1987 -71 1999 -37
rect -2045 -77 -1987 -71
rect -1853 -77 -1795 -71
rect -1661 -77 -1603 -71
rect -1469 -77 -1411 -71
rect -1277 -77 -1219 -71
rect -1085 -77 -1027 -71
rect -893 -77 -835 -71
rect -701 -77 -643 -71
rect -509 -77 -451 -71
rect -317 -77 -259 -71
rect -125 -77 -67 -71
rect 67 -77 125 -71
rect 259 -77 317 -71
rect 451 -77 509 -71
rect 643 -77 701 -71
rect 835 -77 893 -71
rect 1027 -77 1085 -71
rect 1219 -77 1277 -71
rect 1411 -77 1469 -71
rect 1603 -77 1661 -71
rect 1795 -77 1853 -71
rect 1987 -77 2045 -71
rect -2141 -565 -2083 -559
rect -1949 -565 -1891 -559
rect -1757 -565 -1699 -559
rect -1565 -565 -1507 -559
rect -1373 -565 -1315 -559
rect -1181 -565 -1123 -559
rect -989 -565 -931 -559
rect -797 -565 -739 -559
rect -605 -565 -547 -559
rect -413 -565 -355 -559
rect -221 -565 -163 -559
rect -29 -565 29 -559
rect 163 -565 221 -559
rect 355 -565 413 -559
rect 547 -565 605 -559
rect 739 -565 797 -559
rect 931 -565 989 -559
rect 1123 -565 1181 -559
rect 1315 -565 1373 -559
rect 1507 -565 1565 -559
rect 1699 -565 1757 -559
rect 1891 -565 1949 -559
rect 2083 -565 2141 -559
rect -2141 -599 -2129 -565
rect -1949 -599 -1937 -565
rect -1757 -599 -1745 -565
rect -1565 -599 -1553 -565
rect -1373 -599 -1361 -565
rect -1181 -599 -1169 -565
rect -989 -599 -977 -565
rect -797 -599 -785 -565
rect -605 -599 -593 -565
rect -413 -599 -401 -565
rect -221 -599 -209 -565
rect -29 -599 -17 -565
rect 163 -599 175 -565
rect 355 -599 367 -565
rect 547 -599 559 -565
rect 739 -599 751 -565
rect 931 -599 943 -565
rect 1123 -599 1135 -565
rect 1315 -599 1327 -565
rect 1507 -599 1519 -565
rect 1699 -599 1711 -565
rect 1891 -599 1903 -565
rect 2083 -599 2095 -565
rect -2141 -605 -2083 -599
rect -1949 -605 -1891 -599
rect -1757 -605 -1699 -599
rect -1565 -605 -1507 -599
rect -1373 -605 -1315 -599
rect -1181 -605 -1123 -599
rect -989 -605 -931 -599
rect -797 -605 -739 -599
rect -605 -605 -547 -599
rect -413 -605 -355 -599
rect -221 -605 -163 -599
rect -29 -605 29 -599
rect 163 -605 221 -599
rect 355 -605 413 -599
rect 547 -605 605 -599
rect 739 -605 797 -599
rect 931 -605 989 -599
rect 1123 -605 1181 -599
rect 1315 -605 1373 -599
rect 1507 -605 1565 -599
rect 1699 -605 1757 -599
rect 1891 -605 1949 -599
rect 2083 -605 2141 -599
<< nwell >>
rect -2327 -737 2327 737
<< pmos >>
rect -2127 118 -2097 518
rect -2031 118 -2001 518
rect -1935 118 -1905 518
rect -1839 118 -1809 518
rect -1743 118 -1713 518
rect -1647 118 -1617 518
rect -1551 118 -1521 518
rect -1455 118 -1425 518
rect -1359 118 -1329 518
rect -1263 118 -1233 518
rect -1167 118 -1137 518
rect -1071 118 -1041 518
rect -975 118 -945 518
rect -879 118 -849 518
rect -783 118 -753 518
rect -687 118 -657 518
rect -591 118 -561 518
rect -495 118 -465 518
rect -399 118 -369 518
rect -303 118 -273 518
rect -207 118 -177 518
rect -111 118 -81 518
rect -15 118 15 518
rect 81 118 111 518
rect 177 118 207 518
rect 273 118 303 518
rect 369 118 399 518
rect 465 118 495 518
rect 561 118 591 518
rect 657 118 687 518
rect 753 118 783 518
rect 849 118 879 518
rect 945 118 975 518
rect 1041 118 1071 518
rect 1137 118 1167 518
rect 1233 118 1263 518
rect 1329 118 1359 518
rect 1425 118 1455 518
rect 1521 118 1551 518
rect 1617 118 1647 518
rect 1713 118 1743 518
rect 1809 118 1839 518
rect 1905 118 1935 518
rect 2001 118 2031 518
rect 2097 118 2127 518
rect -2127 -518 -2097 -118
rect -2031 -518 -2001 -118
rect -1935 -518 -1905 -118
rect -1839 -518 -1809 -118
rect -1743 -518 -1713 -118
rect -1647 -518 -1617 -118
rect -1551 -518 -1521 -118
rect -1455 -518 -1425 -118
rect -1359 -518 -1329 -118
rect -1263 -518 -1233 -118
rect -1167 -518 -1137 -118
rect -1071 -518 -1041 -118
rect -975 -518 -945 -118
rect -879 -518 -849 -118
rect -783 -518 -753 -118
rect -687 -518 -657 -118
rect -591 -518 -561 -118
rect -495 -518 -465 -118
rect -399 -518 -369 -118
rect -303 -518 -273 -118
rect -207 -518 -177 -118
rect -111 -518 -81 -118
rect -15 -518 15 -118
rect 81 -518 111 -118
rect 177 -518 207 -118
rect 273 -518 303 -118
rect 369 -518 399 -118
rect 465 -518 495 -118
rect 561 -518 591 -118
rect 657 -518 687 -118
rect 753 -518 783 -118
rect 849 -518 879 -118
rect 945 -518 975 -118
rect 1041 -518 1071 -118
rect 1137 -518 1167 -118
rect 1233 -518 1263 -118
rect 1329 -518 1359 -118
rect 1425 -518 1455 -118
rect 1521 -518 1551 -118
rect 1617 -518 1647 -118
rect 1713 -518 1743 -118
rect 1809 -518 1839 -118
rect 1905 -518 1935 -118
rect 2001 -518 2031 -118
rect 2097 -518 2127 -118
<< pdiff >>
rect -2189 506 -2127 518
rect -2189 130 -2177 506
rect -2143 130 -2127 506
rect -2189 118 -2127 130
rect -2097 506 -2031 518
rect -2097 130 -2081 506
rect -2047 130 -2031 506
rect -2097 118 -2031 130
rect -2001 506 -1935 518
rect -2001 130 -1985 506
rect -1951 130 -1935 506
rect -2001 118 -1935 130
rect -1905 506 -1839 518
rect -1905 130 -1889 506
rect -1855 130 -1839 506
rect -1905 118 -1839 130
rect -1809 506 -1743 518
rect -1809 130 -1793 506
rect -1759 130 -1743 506
rect -1809 118 -1743 130
rect -1713 506 -1647 518
rect -1713 130 -1697 506
rect -1663 130 -1647 506
rect -1713 118 -1647 130
rect -1617 506 -1551 518
rect -1617 130 -1601 506
rect -1567 130 -1551 506
rect -1617 118 -1551 130
rect -1521 506 -1455 518
rect -1521 130 -1505 506
rect -1471 130 -1455 506
rect -1521 118 -1455 130
rect -1425 506 -1359 518
rect -1425 130 -1409 506
rect -1375 130 -1359 506
rect -1425 118 -1359 130
rect -1329 506 -1263 518
rect -1329 130 -1313 506
rect -1279 130 -1263 506
rect -1329 118 -1263 130
rect -1233 506 -1167 518
rect -1233 130 -1217 506
rect -1183 130 -1167 506
rect -1233 118 -1167 130
rect -1137 506 -1071 518
rect -1137 130 -1121 506
rect -1087 130 -1071 506
rect -1137 118 -1071 130
rect -1041 506 -975 518
rect -1041 130 -1025 506
rect -991 130 -975 506
rect -1041 118 -975 130
rect -945 506 -879 518
rect -945 130 -929 506
rect -895 130 -879 506
rect -945 118 -879 130
rect -849 506 -783 518
rect -849 130 -833 506
rect -799 130 -783 506
rect -849 118 -783 130
rect -753 506 -687 518
rect -753 130 -737 506
rect -703 130 -687 506
rect -753 118 -687 130
rect -657 506 -591 518
rect -657 130 -641 506
rect -607 130 -591 506
rect -657 118 -591 130
rect -561 506 -495 518
rect -561 130 -545 506
rect -511 130 -495 506
rect -561 118 -495 130
rect -465 506 -399 518
rect -465 130 -449 506
rect -415 130 -399 506
rect -465 118 -399 130
rect -369 506 -303 518
rect -369 130 -353 506
rect -319 130 -303 506
rect -369 118 -303 130
rect -273 506 -207 518
rect -273 130 -257 506
rect -223 130 -207 506
rect -273 118 -207 130
rect -177 506 -111 518
rect -177 130 -161 506
rect -127 130 -111 506
rect -177 118 -111 130
rect -81 506 -15 518
rect -81 130 -65 506
rect -31 130 -15 506
rect -81 118 -15 130
rect 15 506 81 518
rect 15 130 31 506
rect 65 130 81 506
rect 15 118 81 130
rect 111 506 177 518
rect 111 130 127 506
rect 161 130 177 506
rect 111 118 177 130
rect 207 506 273 518
rect 207 130 223 506
rect 257 130 273 506
rect 207 118 273 130
rect 303 506 369 518
rect 303 130 319 506
rect 353 130 369 506
rect 303 118 369 130
rect 399 506 465 518
rect 399 130 415 506
rect 449 130 465 506
rect 399 118 465 130
rect 495 506 561 518
rect 495 130 511 506
rect 545 130 561 506
rect 495 118 561 130
rect 591 506 657 518
rect 591 130 607 506
rect 641 130 657 506
rect 591 118 657 130
rect 687 506 753 518
rect 687 130 703 506
rect 737 130 753 506
rect 687 118 753 130
rect 783 506 849 518
rect 783 130 799 506
rect 833 130 849 506
rect 783 118 849 130
rect 879 506 945 518
rect 879 130 895 506
rect 929 130 945 506
rect 879 118 945 130
rect 975 506 1041 518
rect 975 130 991 506
rect 1025 130 1041 506
rect 975 118 1041 130
rect 1071 506 1137 518
rect 1071 130 1087 506
rect 1121 130 1137 506
rect 1071 118 1137 130
rect 1167 506 1233 518
rect 1167 130 1183 506
rect 1217 130 1233 506
rect 1167 118 1233 130
rect 1263 506 1329 518
rect 1263 130 1279 506
rect 1313 130 1329 506
rect 1263 118 1329 130
rect 1359 506 1425 518
rect 1359 130 1375 506
rect 1409 130 1425 506
rect 1359 118 1425 130
rect 1455 506 1521 518
rect 1455 130 1471 506
rect 1505 130 1521 506
rect 1455 118 1521 130
rect 1551 506 1617 518
rect 1551 130 1567 506
rect 1601 130 1617 506
rect 1551 118 1617 130
rect 1647 506 1713 518
rect 1647 130 1663 506
rect 1697 130 1713 506
rect 1647 118 1713 130
rect 1743 506 1809 518
rect 1743 130 1759 506
rect 1793 130 1809 506
rect 1743 118 1809 130
rect 1839 506 1905 518
rect 1839 130 1855 506
rect 1889 130 1905 506
rect 1839 118 1905 130
rect 1935 506 2001 518
rect 1935 130 1951 506
rect 1985 130 2001 506
rect 1935 118 2001 130
rect 2031 506 2097 518
rect 2031 130 2047 506
rect 2081 130 2097 506
rect 2031 118 2097 130
rect 2127 506 2189 518
rect 2127 130 2143 506
rect 2177 130 2189 506
rect 2127 118 2189 130
rect -2189 -130 -2127 -118
rect -2189 -506 -2177 -130
rect -2143 -506 -2127 -130
rect -2189 -518 -2127 -506
rect -2097 -130 -2031 -118
rect -2097 -506 -2081 -130
rect -2047 -506 -2031 -130
rect -2097 -518 -2031 -506
rect -2001 -130 -1935 -118
rect -2001 -506 -1985 -130
rect -1951 -506 -1935 -130
rect -2001 -518 -1935 -506
rect -1905 -130 -1839 -118
rect -1905 -506 -1889 -130
rect -1855 -506 -1839 -130
rect -1905 -518 -1839 -506
rect -1809 -130 -1743 -118
rect -1809 -506 -1793 -130
rect -1759 -506 -1743 -130
rect -1809 -518 -1743 -506
rect -1713 -130 -1647 -118
rect -1713 -506 -1697 -130
rect -1663 -506 -1647 -130
rect -1713 -518 -1647 -506
rect -1617 -130 -1551 -118
rect -1617 -506 -1601 -130
rect -1567 -506 -1551 -130
rect -1617 -518 -1551 -506
rect -1521 -130 -1455 -118
rect -1521 -506 -1505 -130
rect -1471 -506 -1455 -130
rect -1521 -518 -1455 -506
rect -1425 -130 -1359 -118
rect -1425 -506 -1409 -130
rect -1375 -506 -1359 -130
rect -1425 -518 -1359 -506
rect -1329 -130 -1263 -118
rect -1329 -506 -1313 -130
rect -1279 -506 -1263 -130
rect -1329 -518 -1263 -506
rect -1233 -130 -1167 -118
rect -1233 -506 -1217 -130
rect -1183 -506 -1167 -130
rect -1233 -518 -1167 -506
rect -1137 -130 -1071 -118
rect -1137 -506 -1121 -130
rect -1087 -506 -1071 -130
rect -1137 -518 -1071 -506
rect -1041 -130 -975 -118
rect -1041 -506 -1025 -130
rect -991 -506 -975 -130
rect -1041 -518 -975 -506
rect -945 -130 -879 -118
rect -945 -506 -929 -130
rect -895 -506 -879 -130
rect -945 -518 -879 -506
rect -849 -130 -783 -118
rect -849 -506 -833 -130
rect -799 -506 -783 -130
rect -849 -518 -783 -506
rect -753 -130 -687 -118
rect -753 -506 -737 -130
rect -703 -506 -687 -130
rect -753 -518 -687 -506
rect -657 -130 -591 -118
rect -657 -506 -641 -130
rect -607 -506 -591 -130
rect -657 -518 -591 -506
rect -561 -130 -495 -118
rect -561 -506 -545 -130
rect -511 -506 -495 -130
rect -561 -518 -495 -506
rect -465 -130 -399 -118
rect -465 -506 -449 -130
rect -415 -506 -399 -130
rect -465 -518 -399 -506
rect -369 -130 -303 -118
rect -369 -506 -353 -130
rect -319 -506 -303 -130
rect -369 -518 -303 -506
rect -273 -130 -207 -118
rect -273 -506 -257 -130
rect -223 -506 -207 -130
rect -273 -518 -207 -506
rect -177 -130 -111 -118
rect -177 -506 -161 -130
rect -127 -506 -111 -130
rect -177 -518 -111 -506
rect -81 -130 -15 -118
rect -81 -506 -65 -130
rect -31 -506 -15 -130
rect -81 -518 -15 -506
rect 15 -130 81 -118
rect 15 -506 31 -130
rect 65 -506 81 -130
rect 15 -518 81 -506
rect 111 -130 177 -118
rect 111 -506 127 -130
rect 161 -506 177 -130
rect 111 -518 177 -506
rect 207 -130 273 -118
rect 207 -506 223 -130
rect 257 -506 273 -130
rect 207 -518 273 -506
rect 303 -130 369 -118
rect 303 -506 319 -130
rect 353 -506 369 -130
rect 303 -518 369 -506
rect 399 -130 465 -118
rect 399 -506 415 -130
rect 449 -506 465 -130
rect 399 -518 465 -506
rect 495 -130 561 -118
rect 495 -506 511 -130
rect 545 -506 561 -130
rect 495 -518 561 -506
rect 591 -130 657 -118
rect 591 -506 607 -130
rect 641 -506 657 -130
rect 591 -518 657 -506
rect 687 -130 753 -118
rect 687 -506 703 -130
rect 737 -506 753 -130
rect 687 -518 753 -506
rect 783 -130 849 -118
rect 783 -506 799 -130
rect 833 -506 849 -130
rect 783 -518 849 -506
rect 879 -130 945 -118
rect 879 -506 895 -130
rect 929 -506 945 -130
rect 879 -518 945 -506
rect 975 -130 1041 -118
rect 975 -506 991 -130
rect 1025 -506 1041 -130
rect 975 -518 1041 -506
rect 1071 -130 1137 -118
rect 1071 -506 1087 -130
rect 1121 -506 1137 -130
rect 1071 -518 1137 -506
rect 1167 -130 1233 -118
rect 1167 -506 1183 -130
rect 1217 -506 1233 -130
rect 1167 -518 1233 -506
rect 1263 -130 1329 -118
rect 1263 -506 1279 -130
rect 1313 -506 1329 -130
rect 1263 -518 1329 -506
rect 1359 -130 1425 -118
rect 1359 -506 1375 -130
rect 1409 -506 1425 -130
rect 1359 -518 1425 -506
rect 1455 -130 1521 -118
rect 1455 -506 1471 -130
rect 1505 -506 1521 -130
rect 1455 -518 1521 -506
rect 1551 -130 1617 -118
rect 1551 -506 1567 -130
rect 1601 -506 1617 -130
rect 1551 -518 1617 -506
rect 1647 -130 1713 -118
rect 1647 -506 1663 -130
rect 1697 -506 1713 -130
rect 1647 -518 1713 -506
rect 1743 -130 1809 -118
rect 1743 -506 1759 -130
rect 1793 -506 1809 -130
rect 1743 -518 1809 -506
rect 1839 -130 1905 -118
rect 1839 -506 1855 -130
rect 1889 -506 1905 -130
rect 1839 -518 1905 -506
rect 1935 -130 2001 -118
rect 1935 -506 1951 -130
rect 1985 -506 2001 -130
rect 1935 -518 2001 -506
rect 2031 -130 2097 -118
rect 2031 -506 2047 -130
rect 2081 -506 2097 -130
rect 2031 -518 2097 -506
rect 2127 -130 2189 -118
rect 2127 -506 2143 -130
rect 2177 -506 2189 -130
rect 2127 -518 2189 -506
<< pdiffc >>
rect -2177 130 -2143 506
rect -2081 130 -2047 506
rect -1985 130 -1951 506
rect -1889 130 -1855 506
rect -1793 130 -1759 506
rect -1697 130 -1663 506
rect -1601 130 -1567 506
rect -1505 130 -1471 506
rect -1409 130 -1375 506
rect -1313 130 -1279 506
rect -1217 130 -1183 506
rect -1121 130 -1087 506
rect -1025 130 -991 506
rect -929 130 -895 506
rect -833 130 -799 506
rect -737 130 -703 506
rect -641 130 -607 506
rect -545 130 -511 506
rect -449 130 -415 506
rect -353 130 -319 506
rect -257 130 -223 506
rect -161 130 -127 506
rect -65 130 -31 506
rect 31 130 65 506
rect 127 130 161 506
rect 223 130 257 506
rect 319 130 353 506
rect 415 130 449 506
rect 511 130 545 506
rect 607 130 641 506
rect 703 130 737 506
rect 799 130 833 506
rect 895 130 929 506
rect 991 130 1025 506
rect 1087 130 1121 506
rect 1183 130 1217 506
rect 1279 130 1313 506
rect 1375 130 1409 506
rect 1471 130 1505 506
rect 1567 130 1601 506
rect 1663 130 1697 506
rect 1759 130 1793 506
rect 1855 130 1889 506
rect 1951 130 1985 506
rect 2047 130 2081 506
rect 2143 130 2177 506
rect -2177 -506 -2143 -130
rect -2081 -506 -2047 -130
rect -1985 -506 -1951 -130
rect -1889 -506 -1855 -130
rect -1793 -506 -1759 -130
rect -1697 -506 -1663 -130
rect -1601 -506 -1567 -130
rect -1505 -506 -1471 -130
rect -1409 -506 -1375 -130
rect -1313 -506 -1279 -130
rect -1217 -506 -1183 -130
rect -1121 -506 -1087 -130
rect -1025 -506 -991 -130
rect -929 -506 -895 -130
rect -833 -506 -799 -130
rect -737 -506 -703 -130
rect -641 -506 -607 -130
rect -545 -506 -511 -130
rect -449 -506 -415 -130
rect -353 -506 -319 -130
rect -257 -506 -223 -130
rect -161 -506 -127 -130
rect -65 -506 -31 -130
rect 31 -506 65 -130
rect 127 -506 161 -130
rect 223 -506 257 -130
rect 319 -506 353 -130
rect 415 -506 449 -130
rect 511 -506 545 -130
rect 607 -506 641 -130
rect 703 -506 737 -130
rect 799 -506 833 -130
rect 895 -506 929 -130
rect 991 -506 1025 -130
rect 1087 -506 1121 -130
rect 1183 -506 1217 -130
rect 1279 -506 1313 -130
rect 1375 -506 1409 -130
rect 1471 -506 1505 -130
rect 1567 -506 1601 -130
rect 1663 -506 1697 -130
rect 1759 -506 1793 -130
rect 1855 -506 1889 -130
rect 1951 -506 1985 -130
rect 2047 -506 2081 -130
rect 2143 -506 2177 -130
<< nsubdiff >>
rect -2291 667 -2195 701
rect 2195 667 2291 701
rect -2291 605 -2257 667
rect 2257 605 2291 667
rect -2291 -667 -2257 -605
rect 2257 -667 2291 -605
rect -2291 -701 -2195 -667
rect 2195 -701 2291 -667
<< nsubdiffcont >>
rect -2195 667 2195 701
rect -2291 -605 -2257 605
rect 2257 -605 2291 605
rect -2195 -701 2195 -667
<< poly >>
rect -2145 599 -2079 615
rect -2145 565 -2129 599
rect -2095 565 -2079 599
rect -2145 549 -2079 565
rect -1953 599 -1887 615
rect -1953 565 -1937 599
rect -1903 565 -1887 599
rect -1953 549 -1887 565
rect -1761 599 -1695 615
rect -1761 565 -1745 599
rect -1711 565 -1695 599
rect -1761 549 -1695 565
rect -1569 599 -1503 615
rect -1569 565 -1553 599
rect -1519 565 -1503 599
rect -1569 549 -1503 565
rect -1377 599 -1311 615
rect -1377 565 -1361 599
rect -1327 565 -1311 599
rect -1377 549 -1311 565
rect -1185 599 -1119 615
rect -1185 565 -1169 599
rect -1135 565 -1119 599
rect -1185 549 -1119 565
rect -993 599 -927 615
rect -993 565 -977 599
rect -943 565 -927 599
rect -993 549 -927 565
rect -801 599 -735 615
rect -801 565 -785 599
rect -751 565 -735 599
rect -801 549 -735 565
rect -609 599 -543 615
rect -609 565 -593 599
rect -559 565 -543 599
rect -609 549 -543 565
rect -417 599 -351 615
rect -417 565 -401 599
rect -367 565 -351 599
rect -417 549 -351 565
rect -225 599 -159 615
rect -225 565 -209 599
rect -175 565 -159 599
rect -225 549 -159 565
rect -33 599 33 615
rect -33 565 -17 599
rect 17 565 33 599
rect -33 549 33 565
rect 159 599 225 615
rect 159 565 175 599
rect 209 565 225 599
rect 159 549 225 565
rect 351 599 417 615
rect 351 565 367 599
rect 401 565 417 599
rect 351 549 417 565
rect 543 599 609 615
rect 543 565 559 599
rect 593 565 609 599
rect 543 549 609 565
rect 735 599 801 615
rect 735 565 751 599
rect 785 565 801 599
rect 735 549 801 565
rect 927 599 993 615
rect 927 565 943 599
rect 977 565 993 599
rect 927 549 993 565
rect 1119 599 1185 615
rect 1119 565 1135 599
rect 1169 565 1185 599
rect 1119 549 1185 565
rect 1311 599 1377 615
rect 1311 565 1327 599
rect 1361 565 1377 599
rect 1311 549 1377 565
rect 1503 599 1569 615
rect 1503 565 1519 599
rect 1553 565 1569 599
rect 1503 549 1569 565
rect 1695 599 1761 615
rect 1695 565 1711 599
rect 1745 565 1761 599
rect 1695 549 1761 565
rect 1887 599 1953 615
rect 1887 565 1903 599
rect 1937 565 1953 599
rect 1887 549 1953 565
rect 2079 599 2145 615
rect 2079 565 2095 599
rect 2129 565 2145 599
rect 2079 549 2145 565
rect -2127 518 -2097 549
rect -2031 518 -2001 544
rect -1935 518 -1905 549
rect -1839 518 -1809 544
rect -1743 518 -1713 549
rect -1647 518 -1617 544
rect -1551 518 -1521 549
rect -1455 518 -1425 544
rect -1359 518 -1329 549
rect -1263 518 -1233 544
rect -1167 518 -1137 549
rect -1071 518 -1041 544
rect -975 518 -945 549
rect -879 518 -849 544
rect -783 518 -753 549
rect -687 518 -657 544
rect -591 518 -561 549
rect -495 518 -465 544
rect -399 518 -369 549
rect -303 518 -273 544
rect -207 518 -177 549
rect -111 518 -81 544
rect -15 518 15 549
rect 81 518 111 544
rect 177 518 207 549
rect 273 518 303 544
rect 369 518 399 549
rect 465 518 495 544
rect 561 518 591 549
rect 657 518 687 544
rect 753 518 783 549
rect 849 518 879 544
rect 945 518 975 549
rect 1041 518 1071 544
rect 1137 518 1167 549
rect 1233 518 1263 544
rect 1329 518 1359 549
rect 1425 518 1455 544
rect 1521 518 1551 549
rect 1617 518 1647 544
rect 1713 518 1743 549
rect 1809 518 1839 544
rect 1905 518 1935 549
rect 2001 518 2031 544
rect 2097 518 2127 549
rect -2127 92 -2097 118
rect -2031 87 -2001 118
rect -1935 92 -1905 118
rect -1839 87 -1809 118
rect -1743 92 -1713 118
rect -1647 87 -1617 118
rect -1551 92 -1521 118
rect -1455 87 -1425 118
rect -1359 92 -1329 118
rect -1263 87 -1233 118
rect -1167 92 -1137 118
rect -1071 87 -1041 118
rect -975 92 -945 118
rect -879 87 -849 118
rect -783 92 -753 118
rect -687 87 -657 118
rect -591 92 -561 118
rect -495 87 -465 118
rect -399 92 -369 118
rect -303 87 -273 118
rect -207 92 -177 118
rect -111 87 -81 118
rect -15 92 15 118
rect 81 87 111 118
rect 177 92 207 118
rect 273 87 303 118
rect 369 92 399 118
rect 465 87 495 118
rect 561 92 591 118
rect 657 87 687 118
rect 753 92 783 118
rect 849 87 879 118
rect 945 92 975 118
rect 1041 87 1071 118
rect 1137 92 1167 118
rect 1233 87 1263 118
rect 1329 92 1359 118
rect 1425 87 1455 118
rect 1521 92 1551 118
rect 1617 87 1647 118
rect 1713 92 1743 118
rect 1809 87 1839 118
rect 1905 92 1935 118
rect 2001 87 2031 118
rect 2097 92 2127 118
rect -2049 71 -1983 87
rect -2049 37 -2033 71
rect -1999 37 -1983 71
rect -2049 21 -1983 37
rect -1857 71 -1791 87
rect -1857 37 -1841 71
rect -1807 37 -1791 71
rect -1857 21 -1791 37
rect -1665 71 -1599 87
rect -1665 37 -1649 71
rect -1615 37 -1599 71
rect -1665 21 -1599 37
rect -1473 71 -1407 87
rect -1473 37 -1457 71
rect -1423 37 -1407 71
rect -1473 21 -1407 37
rect -1281 71 -1215 87
rect -1281 37 -1265 71
rect -1231 37 -1215 71
rect -1281 21 -1215 37
rect -1089 71 -1023 87
rect -1089 37 -1073 71
rect -1039 37 -1023 71
rect -1089 21 -1023 37
rect -897 71 -831 87
rect -897 37 -881 71
rect -847 37 -831 71
rect -897 21 -831 37
rect -705 71 -639 87
rect -705 37 -689 71
rect -655 37 -639 71
rect -705 21 -639 37
rect -513 71 -447 87
rect -513 37 -497 71
rect -463 37 -447 71
rect -513 21 -447 37
rect -321 71 -255 87
rect -321 37 -305 71
rect -271 37 -255 71
rect -321 21 -255 37
rect -129 71 -63 87
rect -129 37 -113 71
rect -79 37 -63 71
rect -129 21 -63 37
rect 63 71 129 87
rect 63 37 79 71
rect 113 37 129 71
rect 63 21 129 37
rect 255 71 321 87
rect 255 37 271 71
rect 305 37 321 71
rect 255 21 321 37
rect 447 71 513 87
rect 447 37 463 71
rect 497 37 513 71
rect 447 21 513 37
rect 639 71 705 87
rect 639 37 655 71
rect 689 37 705 71
rect 639 21 705 37
rect 831 71 897 87
rect 831 37 847 71
rect 881 37 897 71
rect 831 21 897 37
rect 1023 71 1089 87
rect 1023 37 1039 71
rect 1073 37 1089 71
rect 1023 21 1089 37
rect 1215 71 1281 87
rect 1215 37 1231 71
rect 1265 37 1281 71
rect 1215 21 1281 37
rect 1407 71 1473 87
rect 1407 37 1423 71
rect 1457 37 1473 71
rect 1407 21 1473 37
rect 1599 71 1665 87
rect 1599 37 1615 71
rect 1649 37 1665 71
rect 1599 21 1665 37
rect 1791 71 1857 87
rect 1791 37 1807 71
rect 1841 37 1857 71
rect 1791 21 1857 37
rect 1983 71 2049 87
rect 1983 37 1999 71
rect 2033 37 2049 71
rect 1983 21 2049 37
rect -2049 -37 -1983 -21
rect -2049 -71 -2033 -37
rect -1999 -71 -1983 -37
rect -2049 -87 -1983 -71
rect -1857 -37 -1791 -21
rect -1857 -71 -1841 -37
rect -1807 -71 -1791 -37
rect -1857 -87 -1791 -71
rect -1665 -37 -1599 -21
rect -1665 -71 -1649 -37
rect -1615 -71 -1599 -37
rect -1665 -87 -1599 -71
rect -1473 -37 -1407 -21
rect -1473 -71 -1457 -37
rect -1423 -71 -1407 -37
rect -1473 -87 -1407 -71
rect -1281 -37 -1215 -21
rect -1281 -71 -1265 -37
rect -1231 -71 -1215 -37
rect -1281 -87 -1215 -71
rect -1089 -37 -1023 -21
rect -1089 -71 -1073 -37
rect -1039 -71 -1023 -37
rect -1089 -87 -1023 -71
rect -897 -37 -831 -21
rect -897 -71 -881 -37
rect -847 -71 -831 -37
rect -897 -87 -831 -71
rect -705 -37 -639 -21
rect -705 -71 -689 -37
rect -655 -71 -639 -37
rect -705 -87 -639 -71
rect -513 -37 -447 -21
rect -513 -71 -497 -37
rect -463 -71 -447 -37
rect -513 -87 -447 -71
rect -321 -37 -255 -21
rect -321 -71 -305 -37
rect -271 -71 -255 -37
rect -321 -87 -255 -71
rect -129 -37 -63 -21
rect -129 -71 -113 -37
rect -79 -71 -63 -37
rect -129 -87 -63 -71
rect 63 -37 129 -21
rect 63 -71 79 -37
rect 113 -71 129 -37
rect 63 -87 129 -71
rect 255 -37 321 -21
rect 255 -71 271 -37
rect 305 -71 321 -37
rect 255 -87 321 -71
rect 447 -37 513 -21
rect 447 -71 463 -37
rect 497 -71 513 -37
rect 447 -87 513 -71
rect 639 -37 705 -21
rect 639 -71 655 -37
rect 689 -71 705 -37
rect 639 -87 705 -71
rect 831 -37 897 -21
rect 831 -71 847 -37
rect 881 -71 897 -37
rect 831 -87 897 -71
rect 1023 -37 1089 -21
rect 1023 -71 1039 -37
rect 1073 -71 1089 -37
rect 1023 -87 1089 -71
rect 1215 -37 1281 -21
rect 1215 -71 1231 -37
rect 1265 -71 1281 -37
rect 1215 -87 1281 -71
rect 1407 -37 1473 -21
rect 1407 -71 1423 -37
rect 1457 -71 1473 -37
rect 1407 -87 1473 -71
rect 1599 -37 1665 -21
rect 1599 -71 1615 -37
rect 1649 -71 1665 -37
rect 1599 -87 1665 -71
rect 1791 -37 1857 -21
rect 1791 -71 1807 -37
rect 1841 -71 1857 -37
rect 1791 -87 1857 -71
rect 1983 -37 2049 -21
rect 1983 -71 1999 -37
rect 2033 -71 2049 -37
rect 1983 -87 2049 -71
rect -2127 -118 -2097 -92
rect -2031 -118 -2001 -87
rect -1935 -118 -1905 -92
rect -1839 -118 -1809 -87
rect -1743 -118 -1713 -92
rect -1647 -118 -1617 -87
rect -1551 -118 -1521 -92
rect -1455 -118 -1425 -87
rect -1359 -118 -1329 -92
rect -1263 -118 -1233 -87
rect -1167 -118 -1137 -92
rect -1071 -118 -1041 -87
rect -975 -118 -945 -92
rect -879 -118 -849 -87
rect -783 -118 -753 -92
rect -687 -118 -657 -87
rect -591 -118 -561 -92
rect -495 -118 -465 -87
rect -399 -118 -369 -92
rect -303 -118 -273 -87
rect -207 -118 -177 -92
rect -111 -118 -81 -87
rect -15 -118 15 -92
rect 81 -118 111 -87
rect 177 -118 207 -92
rect 273 -118 303 -87
rect 369 -118 399 -92
rect 465 -118 495 -87
rect 561 -118 591 -92
rect 657 -118 687 -87
rect 753 -118 783 -92
rect 849 -118 879 -87
rect 945 -118 975 -92
rect 1041 -118 1071 -87
rect 1137 -118 1167 -92
rect 1233 -118 1263 -87
rect 1329 -118 1359 -92
rect 1425 -118 1455 -87
rect 1521 -118 1551 -92
rect 1617 -118 1647 -87
rect 1713 -118 1743 -92
rect 1809 -118 1839 -87
rect 1905 -118 1935 -92
rect 2001 -118 2031 -87
rect 2097 -118 2127 -92
rect -2127 -549 -2097 -518
rect -2031 -544 -2001 -518
rect -1935 -549 -1905 -518
rect -1839 -544 -1809 -518
rect -1743 -549 -1713 -518
rect -1647 -544 -1617 -518
rect -1551 -549 -1521 -518
rect -1455 -544 -1425 -518
rect -1359 -549 -1329 -518
rect -1263 -544 -1233 -518
rect -1167 -549 -1137 -518
rect -1071 -544 -1041 -518
rect -975 -549 -945 -518
rect -879 -544 -849 -518
rect -783 -549 -753 -518
rect -687 -544 -657 -518
rect -591 -549 -561 -518
rect -495 -544 -465 -518
rect -399 -549 -369 -518
rect -303 -544 -273 -518
rect -207 -549 -177 -518
rect -111 -544 -81 -518
rect -15 -549 15 -518
rect 81 -544 111 -518
rect 177 -549 207 -518
rect 273 -544 303 -518
rect 369 -549 399 -518
rect 465 -544 495 -518
rect 561 -549 591 -518
rect 657 -544 687 -518
rect 753 -549 783 -518
rect 849 -544 879 -518
rect 945 -549 975 -518
rect 1041 -544 1071 -518
rect 1137 -549 1167 -518
rect 1233 -544 1263 -518
rect 1329 -549 1359 -518
rect 1425 -544 1455 -518
rect 1521 -549 1551 -518
rect 1617 -544 1647 -518
rect 1713 -549 1743 -518
rect 1809 -544 1839 -518
rect 1905 -549 1935 -518
rect 2001 -544 2031 -518
rect 2097 -549 2127 -518
rect -2145 -565 -2079 -549
rect -2145 -599 -2129 -565
rect -2095 -599 -2079 -565
rect -2145 -615 -2079 -599
rect -1953 -565 -1887 -549
rect -1953 -599 -1937 -565
rect -1903 -599 -1887 -565
rect -1953 -615 -1887 -599
rect -1761 -565 -1695 -549
rect -1761 -599 -1745 -565
rect -1711 -599 -1695 -565
rect -1761 -615 -1695 -599
rect -1569 -565 -1503 -549
rect -1569 -599 -1553 -565
rect -1519 -599 -1503 -565
rect -1569 -615 -1503 -599
rect -1377 -565 -1311 -549
rect -1377 -599 -1361 -565
rect -1327 -599 -1311 -565
rect -1377 -615 -1311 -599
rect -1185 -565 -1119 -549
rect -1185 -599 -1169 -565
rect -1135 -599 -1119 -565
rect -1185 -615 -1119 -599
rect -993 -565 -927 -549
rect -993 -599 -977 -565
rect -943 -599 -927 -565
rect -993 -615 -927 -599
rect -801 -565 -735 -549
rect -801 -599 -785 -565
rect -751 -599 -735 -565
rect -801 -615 -735 -599
rect -609 -565 -543 -549
rect -609 -599 -593 -565
rect -559 -599 -543 -565
rect -609 -615 -543 -599
rect -417 -565 -351 -549
rect -417 -599 -401 -565
rect -367 -599 -351 -565
rect -417 -615 -351 -599
rect -225 -565 -159 -549
rect -225 -599 -209 -565
rect -175 -599 -159 -565
rect -225 -615 -159 -599
rect -33 -565 33 -549
rect -33 -599 -17 -565
rect 17 -599 33 -565
rect -33 -615 33 -599
rect 159 -565 225 -549
rect 159 -599 175 -565
rect 209 -599 225 -565
rect 159 -615 225 -599
rect 351 -565 417 -549
rect 351 -599 367 -565
rect 401 -599 417 -565
rect 351 -615 417 -599
rect 543 -565 609 -549
rect 543 -599 559 -565
rect 593 -599 609 -565
rect 543 -615 609 -599
rect 735 -565 801 -549
rect 735 -599 751 -565
rect 785 -599 801 -565
rect 735 -615 801 -599
rect 927 -565 993 -549
rect 927 -599 943 -565
rect 977 -599 993 -565
rect 927 -615 993 -599
rect 1119 -565 1185 -549
rect 1119 -599 1135 -565
rect 1169 -599 1185 -565
rect 1119 -615 1185 -599
rect 1311 -565 1377 -549
rect 1311 -599 1327 -565
rect 1361 -599 1377 -565
rect 1311 -615 1377 -599
rect 1503 -565 1569 -549
rect 1503 -599 1519 -565
rect 1553 -599 1569 -565
rect 1503 -615 1569 -599
rect 1695 -565 1761 -549
rect 1695 -599 1711 -565
rect 1745 -599 1761 -565
rect 1695 -615 1761 -599
rect 1887 -565 1953 -549
rect 1887 -599 1903 -565
rect 1937 -599 1953 -565
rect 1887 -615 1953 -599
rect 2079 -565 2145 -549
rect 2079 -599 2095 -565
rect 2129 -599 2145 -565
rect 2079 -615 2145 -599
<< polycont >>
rect -2129 565 -2095 599
rect -1937 565 -1903 599
rect -1745 565 -1711 599
rect -1553 565 -1519 599
rect -1361 565 -1327 599
rect -1169 565 -1135 599
rect -977 565 -943 599
rect -785 565 -751 599
rect -593 565 -559 599
rect -401 565 -367 599
rect -209 565 -175 599
rect -17 565 17 599
rect 175 565 209 599
rect 367 565 401 599
rect 559 565 593 599
rect 751 565 785 599
rect 943 565 977 599
rect 1135 565 1169 599
rect 1327 565 1361 599
rect 1519 565 1553 599
rect 1711 565 1745 599
rect 1903 565 1937 599
rect 2095 565 2129 599
rect -2033 37 -1999 71
rect -1841 37 -1807 71
rect -1649 37 -1615 71
rect -1457 37 -1423 71
rect -1265 37 -1231 71
rect -1073 37 -1039 71
rect -881 37 -847 71
rect -689 37 -655 71
rect -497 37 -463 71
rect -305 37 -271 71
rect -113 37 -79 71
rect 79 37 113 71
rect 271 37 305 71
rect 463 37 497 71
rect 655 37 689 71
rect 847 37 881 71
rect 1039 37 1073 71
rect 1231 37 1265 71
rect 1423 37 1457 71
rect 1615 37 1649 71
rect 1807 37 1841 71
rect 1999 37 2033 71
rect -2033 -71 -1999 -37
rect -1841 -71 -1807 -37
rect -1649 -71 -1615 -37
rect -1457 -71 -1423 -37
rect -1265 -71 -1231 -37
rect -1073 -71 -1039 -37
rect -881 -71 -847 -37
rect -689 -71 -655 -37
rect -497 -71 -463 -37
rect -305 -71 -271 -37
rect -113 -71 -79 -37
rect 79 -71 113 -37
rect 271 -71 305 -37
rect 463 -71 497 -37
rect 655 -71 689 -37
rect 847 -71 881 -37
rect 1039 -71 1073 -37
rect 1231 -71 1265 -37
rect 1423 -71 1457 -37
rect 1615 -71 1649 -37
rect 1807 -71 1841 -37
rect 1999 -71 2033 -37
rect -2129 -599 -2095 -565
rect -1937 -599 -1903 -565
rect -1745 -599 -1711 -565
rect -1553 -599 -1519 -565
rect -1361 -599 -1327 -565
rect -1169 -599 -1135 -565
rect -977 -599 -943 -565
rect -785 -599 -751 -565
rect -593 -599 -559 -565
rect -401 -599 -367 -565
rect -209 -599 -175 -565
rect -17 -599 17 -565
rect 175 -599 209 -565
rect 367 -599 401 -565
rect 559 -599 593 -565
rect 751 -599 785 -565
rect 943 -599 977 -565
rect 1135 -599 1169 -565
rect 1327 -599 1361 -565
rect 1519 -599 1553 -565
rect 1711 -599 1745 -565
rect 1903 -599 1937 -565
rect 2095 -599 2129 -565
<< locali >>
rect -2291 667 -2195 701
rect 2195 667 2291 701
rect -2291 605 -2257 667
rect 2257 605 2291 667
rect -2145 565 -2129 599
rect -2095 565 -2079 599
rect -1953 565 -1937 599
rect -1903 565 -1887 599
rect -1761 565 -1745 599
rect -1711 565 -1695 599
rect -1569 565 -1553 599
rect -1519 565 -1503 599
rect -1377 565 -1361 599
rect -1327 565 -1311 599
rect -1185 565 -1169 599
rect -1135 565 -1119 599
rect -993 565 -977 599
rect -943 565 -927 599
rect -801 565 -785 599
rect -751 565 -735 599
rect -609 565 -593 599
rect -559 565 -543 599
rect -417 565 -401 599
rect -367 565 -351 599
rect -225 565 -209 599
rect -175 565 -159 599
rect -33 565 -17 599
rect 17 565 33 599
rect 159 565 175 599
rect 209 565 225 599
rect 351 565 367 599
rect 401 565 417 599
rect 543 565 559 599
rect 593 565 609 599
rect 735 565 751 599
rect 785 565 801 599
rect 927 565 943 599
rect 977 565 993 599
rect 1119 565 1135 599
rect 1169 565 1185 599
rect 1311 565 1327 599
rect 1361 565 1377 599
rect 1503 565 1519 599
rect 1553 565 1569 599
rect 1695 565 1711 599
rect 1745 565 1761 599
rect 1887 565 1903 599
rect 1937 565 1953 599
rect 2079 565 2095 599
rect 2129 565 2145 599
rect -2177 506 -2143 522
rect -2177 114 -2143 130
rect -2081 506 -2047 522
rect -2081 114 -2047 130
rect -1985 506 -1951 522
rect -1985 114 -1951 130
rect -1889 506 -1855 522
rect -1889 114 -1855 130
rect -1793 506 -1759 522
rect -1793 114 -1759 130
rect -1697 506 -1663 522
rect -1697 114 -1663 130
rect -1601 506 -1567 522
rect -1601 114 -1567 130
rect -1505 506 -1471 522
rect -1505 114 -1471 130
rect -1409 506 -1375 522
rect -1409 114 -1375 130
rect -1313 506 -1279 522
rect -1313 114 -1279 130
rect -1217 506 -1183 522
rect -1217 114 -1183 130
rect -1121 506 -1087 522
rect -1121 114 -1087 130
rect -1025 506 -991 522
rect -1025 114 -991 130
rect -929 506 -895 522
rect -929 114 -895 130
rect -833 506 -799 522
rect -833 114 -799 130
rect -737 506 -703 522
rect -737 114 -703 130
rect -641 506 -607 522
rect -641 114 -607 130
rect -545 506 -511 522
rect -545 114 -511 130
rect -449 506 -415 522
rect -449 114 -415 130
rect -353 506 -319 522
rect -353 114 -319 130
rect -257 506 -223 522
rect -257 114 -223 130
rect -161 506 -127 522
rect -161 114 -127 130
rect -65 506 -31 522
rect -65 114 -31 130
rect 31 506 65 522
rect 31 114 65 130
rect 127 506 161 522
rect 127 114 161 130
rect 223 506 257 522
rect 223 114 257 130
rect 319 506 353 522
rect 319 114 353 130
rect 415 506 449 522
rect 415 114 449 130
rect 511 506 545 522
rect 511 114 545 130
rect 607 506 641 522
rect 607 114 641 130
rect 703 506 737 522
rect 703 114 737 130
rect 799 506 833 522
rect 799 114 833 130
rect 895 506 929 522
rect 895 114 929 130
rect 991 506 1025 522
rect 991 114 1025 130
rect 1087 506 1121 522
rect 1087 114 1121 130
rect 1183 506 1217 522
rect 1183 114 1217 130
rect 1279 506 1313 522
rect 1279 114 1313 130
rect 1375 506 1409 522
rect 1375 114 1409 130
rect 1471 506 1505 522
rect 1471 114 1505 130
rect 1567 506 1601 522
rect 1567 114 1601 130
rect 1663 506 1697 522
rect 1663 114 1697 130
rect 1759 506 1793 522
rect 1759 114 1793 130
rect 1855 506 1889 522
rect 1855 114 1889 130
rect 1951 506 1985 522
rect 1951 114 1985 130
rect 2047 506 2081 522
rect 2047 114 2081 130
rect 2143 506 2177 522
rect 2143 114 2177 130
rect -2049 37 -2033 71
rect -1999 37 -1983 71
rect -1857 37 -1841 71
rect -1807 37 -1791 71
rect -1665 37 -1649 71
rect -1615 37 -1599 71
rect -1473 37 -1457 71
rect -1423 37 -1407 71
rect -1281 37 -1265 71
rect -1231 37 -1215 71
rect -1089 37 -1073 71
rect -1039 37 -1023 71
rect -897 37 -881 71
rect -847 37 -831 71
rect -705 37 -689 71
rect -655 37 -639 71
rect -513 37 -497 71
rect -463 37 -447 71
rect -321 37 -305 71
rect -271 37 -255 71
rect -129 37 -113 71
rect -79 37 -63 71
rect 63 37 79 71
rect 113 37 129 71
rect 255 37 271 71
rect 305 37 321 71
rect 447 37 463 71
rect 497 37 513 71
rect 639 37 655 71
rect 689 37 705 71
rect 831 37 847 71
rect 881 37 897 71
rect 1023 37 1039 71
rect 1073 37 1089 71
rect 1215 37 1231 71
rect 1265 37 1281 71
rect 1407 37 1423 71
rect 1457 37 1473 71
rect 1599 37 1615 71
rect 1649 37 1665 71
rect 1791 37 1807 71
rect 1841 37 1857 71
rect 1983 37 1999 71
rect 2033 37 2049 71
rect -2049 -71 -2033 -37
rect -1999 -71 -1983 -37
rect -1857 -71 -1841 -37
rect -1807 -71 -1791 -37
rect -1665 -71 -1649 -37
rect -1615 -71 -1599 -37
rect -1473 -71 -1457 -37
rect -1423 -71 -1407 -37
rect -1281 -71 -1265 -37
rect -1231 -71 -1215 -37
rect -1089 -71 -1073 -37
rect -1039 -71 -1023 -37
rect -897 -71 -881 -37
rect -847 -71 -831 -37
rect -705 -71 -689 -37
rect -655 -71 -639 -37
rect -513 -71 -497 -37
rect -463 -71 -447 -37
rect -321 -71 -305 -37
rect -271 -71 -255 -37
rect -129 -71 -113 -37
rect -79 -71 -63 -37
rect 63 -71 79 -37
rect 113 -71 129 -37
rect 255 -71 271 -37
rect 305 -71 321 -37
rect 447 -71 463 -37
rect 497 -71 513 -37
rect 639 -71 655 -37
rect 689 -71 705 -37
rect 831 -71 847 -37
rect 881 -71 897 -37
rect 1023 -71 1039 -37
rect 1073 -71 1089 -37
rect 1215 -71 1231 -37
rect 1265 -71 1281 -37
rect 1407 -71 1423 -37
rect 1457 -71 1473 -37
rect 1599 -71 1615 -37
rect 1649 -71 1665 -37
rect 1791 -71 1807 -37
rect 1841 -71 1857 -37
rect 1983 -71 1999 -37
rect 2033 -71 2049 -37
rect -2177 -130 -2143 -114
rect -2177 -522 -2143 -506
rect -2081 -130 -2047 -114
rect -2081 -522 -2047 -506
rect -1985 -130 -1951 -114
rect -1985 -522 -1951 -506
rect -1889 -130 -1855 -114
rect -1889 -522 -1855 -506
rect -1793 -130 -1759 -114
rect -1793 -522 -1759 -506
rect -1697 -130 -1663 -114
rect -1697 -522 -1663 -506
rect -1601 -130 -1567 -114
rect -1601 -522 -1567 -506
rect -1505 -130 -1471 -114
rect -1505 -522 -1471 -506
rect -1409 -130 -1375 -114
rect -1409 -522 -1375 -506
rect -1313 -130 -1279 -114
rect -1313 -522 -1279 -506
rect -1217 -130 -1183 -114
rect -1217 -522 -1183 -506
rect -1121 -130 -1087 -114
rect -1121 -522 -1087 -506
rect -1025 -130 -991 -114
rect -1025 -522 -991 -506
rect -929 -130 -895 -114
rect -929 -522 -895 -506
rect -833 -130 -799 -114
rect -833 -522 -799 -506
rect -737 -130 -703 -114
rect -737 -522 -703 -506
rect -641 -130 -607 -114
rect -641 -522 -607 -506
rect -545 -130 -511 -114
rect -545 -522 -511 -506
rect -449 -130 -415 -114
rect -449 -522 -415 -506
rect -353 -130 -319 -114
rect -353 -522 -319 -506
rect -257 -130 -223 -114
rect -257 -522 -223 -506
rect -161 -130 -127 -114
rect -161 -522 -127 -506
rect -65 -130 -31 -114
rect -65 -522 -31 -506
rect 31 -130 65 -114
rect 31 -522 65 -506
rect 127 -130 161 -114
rect 127 -522 161 -506
rect 223 -130 257 -114
rect 223 -522 257 -506
rect 319 -130 353 -114
rect 319 -522 353 -506
rect 415 -130 449 -114
rect 415 -522 449 -506
rect 511 -130 545 -114
rect 511 -522 545 -506
rect 607 -130 641 -114
rect 607 -522 641 -506
rect 703 -130 737 -114
rect 703 -522 737 -506
rect 799 -130 833 -114
rect 799 -522 833 -506
rect 895 -130 929 -114
rect 895 -522 929 -506
rect 991 -130 1025 -114
rect 991 -522 1025 -506
rect 1087 -130 1121 -114
rect 1087 -522 1121 -506
rect 1183 -130 1217 -114
rect 1183 -522 1217 -506
rect 1279 -130 1313 -114
rect 1279 -522 1313 -506
rect 1375 -130 1409 -114
rect 1375 -522 1409 -506
rect 1471 -130 1505 -114
rect 1471 -522 1505 -506
rect 1567 -130 1601 -114
rect 1567 -522 1601 -506
rect 1663 -130 1697 -114
rect 1663 -522 1697 -506
rect 1759 -130 1793 -114
rect 1759 -522 1793 -506
rect 1855 -130 1889 -114
rect 1855 -522 1889 -506
rect 1951 -130 1985 -114
rect 1951 -522 1985 -506
rect 2047 -130 2081 -114
rect 2047 -522 2081 -506
rect 2143 -130 2177 -114
rect 2143 -522 2177 -506
rect -2145 -599 -2129 -565
rect -2095 -599 -2079 -565
rect -1953 -599 -1937 -565
rect -1903 -599 -1887 -565
rect -1761 -599 -1745 -565
rect -1711 -599 -1695 -565
rect -1569 -599 -1553 -565
rect -1519 -599 -1503 -565
rect -1377 -599 -1361 -565
rect -1327 -599 -1311 -565
rect -1185 -599 -1169 -565
rect -1135 -599 -1119 -565
rect -993 -599 -977 -565
rect -943 -599 -927 -565
rect -801 -599 -785 -565
rect -751 -599 -735 -565
rect -609 -599 -593 -565
rect -559 -599 -543 -565
rect -417 -599 -401 -565
rect -367 -599 -351 -565
rect -225 -599 -209 -565
rect -175 -599 -159 -565
rect -33 -599 -17 -565
rect 17 -599 33 -565
rect 159 -599 175 -565
rect 209 -599 225 -565
rect 351 -599 367 -565
rect 401 -599 417 -565
rect 543 -599 559 -565
rect 593 -599 609 -565
rect 735 -599 751 -565
rect 785 -599 801 -565
rect 927 -599 943 -565
rect 977 -599 993 -565
rect 1119 -599 1135 -565
rect 1169 -599 1185 -565
rect 1311 -599 1327 -565
rect 1361 -599 1377 -565
rect 1503 -599 1519 -565
rect 1553 -599 1569 -565
rect 1695 -599 1711 -565
rect 1745 -599 1761 -565
rect 1887 -599 1903 -565
rect 1937 -599 1953 -565
rect 2079 -599 2095 -565
rect 2129 -599 2145 -565
rect -2291 -667 -2257 -605
rect 2257 -667 2291 -605
rect -2291 -701 -2195 -667
rect 2195 -701 2291 -667
<< viali >>
rect -2129 565 -2095 599
rect -1937 565 -1903 599
rect -1745 565 -1711 599
rect -1553 565 -1519 599
rect -1361 565 -1327 599
rect -1169 565 -1135 599
rect -977 565 -943 599
rect -785 565 -751 599
rect -593 565 -559 599
rect -401 565 -367 599
rect -209 565 -175 599
rect -17 565 17 599
rect 175 565 209 599
rect 367 565 401 599
rect 559 565 593 599
rect 751 565 785 599
rect 943 565 977 599
rect 1135 565 1169 599
rect 1327 565 1361 599
rect 1519 565 1553 599
rect 1711 565 1745 599
rect 1903 565 1937 599
rect 2095 565 2129 599
rect -2177 130 -2143 506
rect -2081 130 -2047 506
rect -1985 130 -1951 506
rect -1889 130 -1855 506
rect -1793 130 -1759 506
rect -1697 130 -1663 506
rect -1601 130 -1567 506
rect -1505 130 -1471 506
rect -1409 130 -1375 506
rect -1313 130 -1279 506
rect -1217 130 -1183 506
rect -1121 130 -1087 506
rect -1025 130 -991 506
rect -929 130 -895 506
rect -833 130 -799 506
rect -737 130 -703 506
rect -641 130 -607 506
rect -545 130 -511 506
rect -449 130 -415 506
rect -353 130 -319 506
rect -257 130 -223 506
rect -161 130 -127 506
rect -65 130 -31 506
rect 31 130 65 506
rect 127 130 161 506
rect 223 130 257 506
rect 319 130 353 506
rect 415 130 449 506
rect 511 130 545 506
rect 607 130 641 506
rect 703 130 737 506
rect 799 130 833 506
rect 895 130 929 506
rect 991 130 1025 506
rect 1087 130 1121 506
rect 1183 130 1217 506
rect 1279 130 1313 506
rect 1375 130 1409 506
rect 1471 130 1505 506
rect 1567 130 1601 506
rect 1663 130 1697 506
rect 1759 130 1793 506
rect 1855 130 1889 506
rect 1951 130 1985 506
rect 2047 130 2081 506
rect 2143 130 2177 506
rect -2033 37 -1999 71
rect -1841 37 -1807 71
rect -1649 37 -1615 71
rect -1457 37 -1423 71
rect -1265 37 -1231 71
rect -1073 37 -1039 71
rect -881 37 -847 71
rect -689 37 -655 71
rect -497 37 -463 71
rect -305 37 -271 71
rect -113 37 -79 71
rect 79 37 113 71
rect 271 37 305 71
rect 463 37 497 71
rect 655 37 689 71
rect 847 37 881 71
rect 1039 37 1073 71
rect 1231 37 1265 71
rect 1423 37 1457 71
rect 1615 37 1649 71
rect 1807 37 1841 71
rect 1999 37 2033 71
rect -2033 -71 -1999 -37
rect -1841 -71 -1807 -37
rect -1649 -71 -1615 -37
rect -1457 -71 -1423 -37
rect -1265 -71 -1231 -37
rect -1073 -71 -1039 -37
rect -881 -71 -847 -37
rect -689 -71 -655 -37
rect -497 -71 -463 -37
rect -305 -71 -271 -37
rect -113 -71 -79 -37
rect 79 -71 113 -37
rect 271 -71 305 -37
rect 463 -71 497 -37
rect 655 -71 689 -37
rect 847 -71 881 -37
rect 1039 -71 1073 -37
rect 1231 -71 1265 -37
rect 1423 -71 1457 -37
rect 1615 -71 1649 -37
rect 1807 -71 1841 -37
rect 1999 -71 2033 -37
rect -2177 -506 -2143 -130
rect -2081 -506 -2047 -130
rect -1985 -506 -1951 -130
rect -1889 -506 -1855 -130
rect -1793 -506 -1759 -130
rect -1697 -506 -1663 -130
rect -1601 -506 -1567 -130
rect -1505 -506 -1471 -130
rect -1409 -506 -1375 -130
rect -1313 -506 -1279 -130
rect -1217 -506 -1183 -130
rect -1121 -506 -1087 -130
rect -1025 -506 -991 -130
rect -929 -506 -895 -130
rect -833 -506 -799 -130
rect -737 -506 -703 -130
rect -641 -506 -607 -130
rect -545 -506 -511 -130
rect -449 -506 -415 -130
rect -353 -506 -319 -130
rect -257 -506 -223 -130
rect -161 -506 -127 -130
rect -65 -506 -31 -130
rect 31 -506 65 -130
rect 127 -506 161 -130
rect 223 -506 257 -130
rect 319 -506 353 -130
rect 415 -506 449 -130
rect 511 -506 545 -130
rect 607 -506 641 -130
rect 703 -506 737 -130
rect 799 -506 833 -130
rect 895 -506 929 -130
rect 991 -506 1025 -130
rect 1087 -506 1121 -130
rect 1183 -506 1217 -130
rect 1279 -506 1313 -130
rect 1375 -506 1409 -130
rect 1471 -506 1505 -130
rect 1567 -506 1601 -130
rect 1663 -506 1697 -130
rect 1759 -506 1793 -130
rect 1855 -506 1889 -130
rect 1951 -506 1985 -130
rect 2047 -506 2081 -130
rect 2143 -506 2177 -130
rect -2129 -599 -2095 -565
rect -1937 -599 -1903 -565
rect -1745 -599 -1711 -565
rect -1553 -599 -1519 -565
rect -1361 -599 -1327 -565
rect -1169 -599 -1135 -565
rect -977 -599 -943 -565
rect -785 -599 -751 -565
rect -593 -599 -559 -565
rect -401 -599 -367 -565
rect -209 -599 -175 -565
rect -17 -599 17 -565
rect 175 -599 209 -565
rect 367 -599 401 -565
rect 559 -599 593 -565
rect 751 -599 785 -565
rect 943 -599 977 -565
rect 1135 -599 1169 -565
rect 1327 -599 1361 -565
rect 1519 -599 1553 -565
rect 1711 -599 1745 -565
rect 1903 -599 1937 -565
rect 2095 -599 2129 -565
<< metal1 >>
rect -2141 599 -2083 605
rect -2141 565 -2129 599
rect -2095 565 -2083 599
rect -2141 559 -2083 565
rect -1949 599 -1891 605
rect -1949 565 -1937 599
rect -1903 565 -1891 599
rect -1949 559 -1891 565
rect -1757 599 -1699 605
rect -1757 565 -1745 599
rect -1711 565 -1699 599
rect -1757 559 -1699 565
rect -1565 599 -1507 605
rect -1565 565 -1553 599
rect -1519 565 -1507 599
rect -1565 559 -1507 565
rect -1373 599 -1315 605
rect -1373 565 -1361 599
rect -1327 565 -1315 599
rect -1373 559 -1315 565
rect -1181 599 -1123 605
rect -1181 565 -1169 599
rect -1135 565 -1123 599
rect -1181 559 -1123 565
rect -989 599 -931 605
rect -989 565 -977 599
rect -943 565 -931 599
rect -989 559 -931 565
rect -797 599 -739 605
rect -797 565 -785 599
rect -751 565 -739 599
rect -797 559 -739 565
rect -605 599 -547 605
rect -605 565 -593 599
rect -559 565 -547 599
rect -605 559 -547 565
rect -413 599 -355 605
rect -413 565 -401 599
rect -367 565 -355 599
rect -413 559 -355 565
rect -221 599 -163 605
rect -221 565 -209 599
rect -175 565 -163 599
rect -221 559 -163 565
rect -29 599 29 605
rect -29 565 -17 599
rect 17 565 29 599
rect -29 559 29 565
rect 163 599 221 605
rect 163 565 175 599
rect 209 565 221 599
rect 163 559 221 565
rect 355 599 413 605
rect 355 565 367 599
rect 401 565 413 599
rect 355 559 413 565
rect 547 599 605 605
rect 547 565 559 599
rect 593 565 605 599
rect 547 559 605 565
rect 739 599 797 605
rect 739 565 751 599
rect 785 565 797 599
rect 739 559 797 565
rect 931 599 989 605
rect 931 565 943 599
rect 977 565 989 599
rect 931 559 989 565
rect 1123 599 1181 605
rect 1123 565 1135 599
rect 1169 565 1181 599
rect 1123 559 1181 565
rect 1315 599 1373 605
rect 1315 565 1327 599
rect 1361 565 1373 599
rect 1315 559 1373 565
rect 1507 599 1565 605
rect 1507 565 1519 599
rect 1553 565 1565 599
rect 1507 559 1565 565
rect 1699 599 1757 605
rect 1699 565 1711 599
rect 1745 565 1757 599
rect 1699 559 1757 565
rect 1891 599 1949 605
rect 1891 565 1903 599
rect 1937 565 1949 599
rect 1891 559 1949 565
rect 2083 599 2141 605
rect 2083 565 2095 599
rect 2129 565 2141 599
rect 2083 559 2141 565
rect -2183 506 -2137 518
rect -2183 130 -2177 506
rect -2143 130 -2137 506
rect -2183 118 -2137 130
rect -2087 506 -2041 518
rect -2087 130 -2081 506
rect -2047 130 -2041 506
rect -2087 118 -2041 130
rect -1991 506 -1945 518
rect -1991 130 -1985 506
rect -1951 130 -1945 506
rect -1991 118 -1945 130
rect -1895 506 -1849 518
rect -1895 130 -1889 506
rect -1855 130 -1849 506
rect -1895 118 -1849 130
rect -1799 506 -1753 518
rect -1799 130 -1793 506
rect -1759 130 -1753 506
rect -1799 118 -1753 130
rect -1703 506 -1657 518
rect -1703 130 -1697 506
rect -1663 130 -1657 506
rect -1703 118 -1657 130
rect -1607 506 -1561 518
rect -1607 130 -1601 506
rect -1567 130 -1561 506
rect -1607 118 -1561 130
rect -1511 506 -1465 518
rect -1511 130 -1505 506
rect -1471 130 -1465 506
rect -1511 118 -1465 130
rect -1415 506 -1369 518
rect -1415 130 -1409 506
rect -1375 130 -1369 506
rect -1415 118 -1369 130
rect -1319 506 -1273 518
rect -1319 130 -1313 506
rect -1279 130 -1273 506
rect -1319 118 -1273 130
rect -1223 506 -1177 518
rect -1223 130 -1217 506
rect -1183 130 -1177 506
rect -1223 118 -1177 130
rect -1127 506 -1081 518
rect -1127 130 -1121 506
rect -1087 130 -1081 506
rect -1127 118 -1081 130
rect -1031 506 -985 518
rect -1031 130 -1025 506
rect -991 130 -985 506
rect -1031 118 -985 130
rect -935 506 -889 518
rect -935 130 -929 506
rect -895 130 -889 506
rect -935 118 -889 130
rect -839 506 -793 518
rect -839 130 -833 506
rect -799 130 -793 506
rect -839 118 -793 130
rect -743 506 -697 518
rect -743 130 -737 506
rect -703 130 -697 506
rect -743 118 -697 130
rect -647 506 -601 518
rect -647 130 -641 506
rect -607 130 -601 506
rect -647 118 -601 130
rect -551 506 -505 518
rect -551 130 -545 506
rect -511 130 -505 506
rect -551 118 -505 130
rect -455 506 -409 518
rect -455 130 -449 506
rect -415 130 -409 506
rect -455 118 -409 130
rect -359 506 -313 518
rect -359 130 -353 506
rect -319 130 -313 506
rect -359 118 -313 130
rect -263 506 -217 518
rect -263 130 -257 506
rect -223 130 -217 506
rect -263 118 -217 130
rect -167 506 -121 518
rect -167 130 -161 506
rect -127 130 -121 506
rect -167 118 -121 130
rect -71 506 -25 518
rect -71 130 -65 506
rect -31 130 -25 506
rect -71 118 -25 130
rect 25 506 71 518
rect 25 130 31 506
rect 65 130 71 506
rect 25 118 71 130
rect 121 506 167 518
rect 121 130 127 506
rect 161 130 167 506
rect 121 118 167 130
rect 217 506 263 518
rect 217 130 223 506
rect 257 130 263 506
rect 217 118 263 130
rect 313 506 359 518
rect 313 130 319 506
rect 353 130 359 506
rect 313 118 359 130
rect 409 506 455 518
rect 409 130 415 506
rect 449 130 455 506
rect 409 118 455 130
rect 505 506 551 518
rect 505 130 511 506
rect 545 130 551 506
rect 505 118 551 130
rect 601 506 647 518
rect 601 130 607 506
rect 641 130 647 506
rect 601 118 647 130
rect 697 506 743 518
rect 697 130 703 506
rect 737 130 743 506
rect 697 118 743 130
rect 793 506 839 518
rect 793 130 799 506
rect 833 130 839 506
rect 793 118 839 130
rect 889 506 935 518
rect 889 130 895 506
rect 929 130 935 506
rect 889 118 935 130
rect 985 506 1031 518
rect 985 130 991 506
rect 1025 130 1031 506
rect 985 118 1031 130
rect 1081 506 1127 518
rect 1081 130 1087 506
rect 1121 130 1127 506
rect 1081 118 1127 130
rect 1177 506 1223 518
rect 1177 130 1183 506
rect 1217 130 1223 506
rect 1177 118 1223 130
rect 1273 506 1319 518
rect 1273 130 1279 506
rect 1313 130 1319 506
rect 1273 118 1319 130
rect 1369 506 1415 518
rect 1369 130 1375 506
rect 1409 130 1415 506
rect 1369 118 1415 130
rect 1465 506 1511 518
rect 1465 130 1471 506
rect 1505 130 1511 506
rect 1465 118 1511 130
rect 1561 506 1607 518
rect 1561 130 1567 506
rect 1601 130 1607 506
rect 1561 118 1607 130
rect 1657 506 1703 518
rect 1657 130 1663 506
rect 1697 130 1703 506
rect 1657 118 1703 130
rect 1753 506 1799 518
rect 1753 130 1759 506
rect 1793 130 1799 506
rect 1753 118 1799 130
rect 1849 506 1895 518
rect 1849 130 1855 506
rect 1889 130 1895 506
rect 1849 118 1895 130
rect 1945 506 1991 518
rect 1945 130 1951 506
rect 1985 130 1991 506
rect 1945 118 1991 130
rect 2041 506 2087 518
rect 2041 130 2047 506
rect 2081 130 2087 506
rect 2041 118 2087 130
rect 2137 506 2183 518
rect 2137 130 2143 506
rect 2177 130 2183 506
rect 2137 118 2183 130
rect -2045 71 -1987 77
rect -2045 37 -2033 71
rect -1999 37 -1987 71
rect -2045 31 -1987 37
rect -1853 71 -1795 77
rect -1853 37 -1841 71
rect -1807 37 -1795 71
rect -1853 31 -1795 37
rect -1661 71 -1603 77
rect -1661 37 -1649 71
rect -1615 37 -1603 71
rect -1661 31 -1603 37
rect -1469 71 -1411 77
rect -1469 37 -1457 71
rect -1423 37 -1411 71
rect -1469 31 -1411 37
rect -1277 71 -1219 77
rect -1277 37 -1265 71
rect -1231 37 -1219 71
rect -1277 31 -1219 37
rect -1085 71 -1027 77
rect -1085 37 -1073 71
rect -1039 37 -1027 71
rect -1085 31 -1027 37
rect -893 71 -835 77
rect -893 37 -881 71
rect -847 37 -835 71
rect -893 31 -835 37
rect -701 71 -643 77
rect -701 37 -689 71
rect -655 37 -643 71
rect -701 31 -643 37
rect -509 71 -451 77
rect -509 37 -497 71
rect -463 37 -451 71
rect -509 31 -451 37
rect -317 71 -259 77
rect -317 37 -305 71
rect -271 37 -259 71
rect -317 31 -259 37
rect -125 71 -67 77
rect -125 37 -113 71
rect -79 37 -67 71
rect -125 31 -67 37
rect 67 71 125 77
rect 67 37 79 71
rect 113 37 125 71
rect 67 31 125 37
rect 259 71 317 77
rect 259 37 271 71
rect 305 37 317 71
rect 259 31 317 37
rect 451 71 509 77
rect 451 37 463 71
rect 497 37 509 71
rect 451 31 509 37
rect 643 71 701 77
rect 643 37 655 71
rect 689 37 701 71
rect 643 31 701 37
rect 835 71 893 77
rect 835 37 847 71
rect 881 37 893 71
rect 835 31 893 37
rect 1027 71 1085 77
rect 1027 37 1039 71
rect 1073 37 1085 71
rect 1027 31 1085 37
rect 1219 71 1277 77
rect 1219 37 1231 71
rect 1265 37 1277 71
rect 1219 31 1277 37
rect 1411 71 1469 77
rect 1411 37 1423 71
rect 1457 37 1469 71
rect 1411 31 1469 37
rect 1603 71 1661 77
rect 1603 37 1615 71
rect 1649 37 1661 71
rect 1603 31 1661 37
rect 1795 71 1853 77
rect 1795 37 1807 71
rect 1841 37 1853 71
rect 1795 31 1853 37
rect 1987 71 2045 77
rect 1987 37 1999 71
rect 2033 37 2045 71
rect 1987 31 2045 37
rect -2045 -37 -1987 -31
rect -2045 -71 -2033 -37
rect -1999 -71 -1987 -37
rect -2045 -77 -1987 -71
rect -1853 -37 -1795 -31
rect -1853 -71 -1841 -37
rect -1807 -71 -1795 -37
rect -1853 -77 -1795 -71
rect -1661 -37 -1603 -31
rect -1661 -71 -1649 -37
rect -1615 -71 -1603 -37
rect -1661 -77 -1603 -71
rect -1469 -37 -1411 -31
rect -1469 -71 -1457 -37
rect -1423 -71 -1411 -37
rect -1469 -77 -1411 -71
rect -1277 -37 -1219 -31
rect -1277 -71 -1265 -37
rect -1231 -71 -1219 -37
rect -1277 -77 -1219 -71
rect -1085 -37 -1027 -31
rect -1085 -71 -1073 -37
rect -1039 -71 -1027 -37
rect -1085 -77 -1027 -71
rect -893 -37 -835 -31
rect -893 -71 -881 -37
rect -847 -71 -835 -37
rect -893 -77 -835 -71
rect -701 -37 -643 -31
rect -701 -71 -689 -37
rect -655 -71 -643 -37
rect -701 -77 -643 -71
rect -509 -37 -451 -31
rect -509 -71 -497 -37
rect -463 -71 -451 -37
rect -509 -77 -451 -71
rect -317 -37 -259 -31
rect -317 -71 -305 -37
rect -271 -71 -259 -37
rect -317 -77 -259 -71
rect -125 -37 -67 -31
rect -125 -71 -113 -37
rect -79 -71 -67 -37
rect -125 -77 -67 -71
rect 67 -37 125 -31
rect 67 -71 79 -37
rect 113 -71 125 -37
rect 67 -77 125 -71
rect 259 -37 317 -31
rect 259 -71 271 -37
rect 305 -71 317 -37
rect 259 -77 317 -71
rect 451 -37 509 -31
rect 451 -71 463 -37
rect 497 -71 509 -37
rect 451 -77 509 -71
rect 643 -37 701 -31
rect 643 -71 655 -37
rect 689 -71 701 -37
rect 643 -77 701 -71
rect 835 -37 893 -31
rect 835 -71 847 -37
rect 881 -71 893 -37
rect 835 -77 893 -71
rect 1027 -37 1085 -31
rect 1027 -71 1039 -37
rect 1073 -71 1085 -37
rect 1027 -77 1085 -71
rect 1219 -37 1277 -31
rect 1219 -71 1231 -37
rect 1265 -71 1277 -37
rect 1219 -77 1277 -71
rect 1411 -37 1469 -31
rect 1411 -71 1423 -37
rect 1457 -71 1469 -37
rect 1411 -77 1469 -71
rect 1603 -37 1661 -31
rect 1603 -71 1615 -37
rect 1649 -71 1661 -37
rect 1603 -77 1661 -71
rect 1795 -37 1853 -31
rect 1795 -71 1807 -37
rect 1841 -71 1853 -37
rect 1795 -77 1853 -71
rect 1987 -37 2045 -31
rect 1987 -71 1999 -37
rect 2033 -71 2045 -37
rect 1987 -77 2045 -71
rect -2183 -130 -2137 -118
rect -2183 -506 -2177 -130
rect -2143 -506 -2137 -130
rect -2183 -518 -2137 -506
rect -2087 -130 -2041 -118
rect -2087 -506 -2081 -130
rect -2047 -506 -2041 -130
rect -2087 -518 -2041 -506
rect -1991 -130 -1945 -118
rect -1991 -506 -1985 -130
rect -1951 -506 -1945 -130
rect -1991 -518 -1945 -506
rect -1895 -130 -1849 -118
rect -1895 -506 -1889 -130
rect -1855 -506 -1849 -130
rect -1895 -518 -1849 -506
rect -1799 -130 -1753 -118
rect -1799 -506 -1793 -130
rect -1759 -506 -1753 -130
rect -1799 -518 -1753 -506
rect -1703 -130 -1657 -118
rect -1703 -506 -1697 -130
rect -1663 -506 -1657 -130
rect -1703 -518 -1657 -506
rect -1607 -130 -1561 -118
rect -1607 -506 -1601 -130
rect -1567 -506 -1561 -130
rect -1607 -518 -1561 -506
rect -1511 -130 -1465 -118
rect -1511 -506 -1505 -130
rect -1471 -506 -1465 -130
rect -1511 -518 -1465 -506
rect -1415 -130 -1369 -118
rect -1415 -506 -1409 -130
rect -1375 -506 -1369 -130
rect -1415 -518 -1369 -506
rect -1319 -130 -1273 -118
rect -1319 -506 -1313 -130
rect -1279 -506 -1273 -130
rect -1319 -518 -1273 -506
rect -1223 -130 -1177 -118
rect -1223 -506 -1217 -130
rect -1183 -506 -1177 -130
rect -1223 -518 -1177 -506
rect -1127 -130 -1081 -118
rect -1127 -506 -1121 -130
rect -1087 -506 -1081 -130
rect -1127 -518 -1081 -506
rect -1031 -130 -985 -118
rect -1031 -506 -1025 -130
rect -991 -506 -985 -130
rect -1031 -518 -985 -506
rect -935 -130 -889 -118
rect -935 -506 -929 -130
rect -895 -506 -889 -130
rect -935 -518 -889 -506
rect -839 -130 -793 -118
rect -839 -506 -833 -130
rect -799 -506 -793 -130
rect -839 -518 -793 -506
rect -743 -130 -697 -118
rect -743 -506 -737 -130
rect -703 -506 -697 -130
rect -743 -518 -697 -506
rect -647 -130 -601 -118
rect -647 -506 -641 -130
rect -607 -506 -601 -130
rect -647 -518 -601 -506
rect -551 -130 -505 -118
rect -551 -506 -545 -130
rect -511 -506 -505 -130
rect -551 -518 -505 -506
rect -455 -130 -409 -118
rect -455 -506 -449 -130
rect -415 -506 -409 -130
rect -455 -518 -409 -506
rect -359 -130 -313 -118
rect -359 -506 -353 -130
rect -319 -506 -313 -130
rect -359 -518 -313 -506
rect -263 -130 -217 -118
rect -263 -506 -257 -130
rect -223 -506 -217 -130
rect -263 -518 -217 -506
rect -167 -130 -121 -118
rect -167 -506 -161 -130
rect -127 -506 -121 -130
rect -167 -518 -121 -506
rect -71 -130 -25 -118
rect -71 -506 -65 -130
rect -31 -506 -25 -130
rect -71 -518 -25 -506
rect 25 -130 71 -118
rect 25 -506 31 -130
rect 65 -506 71 -130
rect 25 -518 71 -506
rect 121 -130 167 -118
rect 121 -506 127 -130
rect 161 -506 167 -130
rect 121 -518 167 -506
rect 217 -130 263 -118
rect 217 -506 223 -130
rect 257 -506 263 -130
rect 217 -518 263 -506
rect 313 -130 359 -118
rect 313 -506 319 -130
rect 353 -506 359 -130
rect 313 -518 359 -506
rect 409 -130 455 -118
rect 409 -506 415 -130
rect 449 -506 455 -130
rect 409 -518 455 -506
rect 505 -130 551 -118
rect 505 -506 511 -130
rect 545 -506 551 -130
rect 505 -518 551 -506
rect 601 -130 647 -118
rect 601 -506 607 -130
rect 641 -506 647 -130
rect 601 -518 647 -506
rect 697 -130 743 -118
rect 697 -506 703 -130
rect 737 -506 743 -130
rect 697 -518 743 -506
rect 793 -130 839 -118
rect 793 -506 799 -130
rect 833 -506 839 -130
rect 793 -518 839 -506
rect 889 -130 935 -118
rect 889 -506 895 -130
rect 929 -506 935 -130
rect 889 -518 935 -506
rect 985 -130 1031 -118
rect 985 -506 991 -130
rect 1025 -506 1031 -130
rect 985 -518 1031 -506
rect 1081 -130 1127 -118
rect 1081 -506 1087 -130
rect 1121 -506 1127 -130
rect 1081 -518 1127 -506
rect 1177 -130 1223 -118
rect 1177 -506 1183 -130
rect 1217 -506 1223 -130
rect 1177 -518 1223 -506
rect 1273 -130 1319 -118
rect 1273 -506 1279 -130
rect 1313 -506 1319 -130
rect 1273 -518 1319 -506
rect 1369 -130 1415 -118
rect 1369 -506 1375 -130
rect 1409 -506 1415 -130
rect 1369 -518 1415 -506
rect 1465 -130 1511 -118
rect 1465 -506 1471 -130
rect 1505 -506 1511 -130
rect 1465 -518 1511 -506
rect 1561 -130 1607 -118
rect 1561 -506 1567 -130
rect 1601 -506 1607 -130
rect 1561 -518 1607 -506
rect 1657 -130 1703 -118
rect 1657 -506 1663 -130
rect 1697 -506 1703 -130
rect 1657 -518 1703 -506
rect 1753 -130 1799 -118
rect 1753 -506 1759 -130
rect 1793 -506 1799 -130
rect 1753 -518 1799 -506
rect 1849 -130 1895 -118
rect 1849 -506 1855 -130
rect 1889 -506 1895 -130
rect 1849 -518 1895 -506
rect 1945 -130 1991 -118
rect 1945 -506 1951 -130
rect 1985 -506 1991 -130
rect 1945 -518 1991 -506
rect 2041 -130 2087 -118
rect 2041 -506 2047 -130
rect 2081 -506 2087 -130
rect 2041 -518 2087 -506
rect 2137 -130 2183 -118
rect 2137 -506 2143 -130
rect 2177 -506 2183 -130
rect 2137 -518 2183 -506
rect -2141 -565 -2083 -559
rect -2141 -599 -2129 -565
rect -2095 -599 -2083 -565
rect -2141 -605 -2083 -599
rect -1949 -565 -1891 -559
rect -1949 -599 -1937 -565
rect -1903 -599 -1891 -565
rect -1949 -605 -1891 -599
rect -1757 -565 -1699 -559
rect -1757 -599 -1745 -565
rect -1711 -599 -1699 -565
rect -1757 -605 -1699 -599
rect -1565 -565 -1507 -559
rect -1565 -599 -1553 -565
rect -1519 -599 -1507 -565
rect -1565 -605 -1507 -599
rect -1373 -565 -1315 -559
rect -1373 -599 -1361 -565
rect -1327 -599 -1315 -565
rect -1373 -605 -1315 -599
rect -1181 -565 -1123 -559
rect -1181 -599 -1169 -565
rect -1135 -599 -1123 -565
rect -1181 -605 -1123 -599
rect -989 -565 -931 -559
rect -989 -599 -977 -565
rect -943 -599 -931 -565
rect -989 -605 -931 -599
rect -797 -565 -739 -559
rect -797 -599 -785 -565
rect -751 -599 -739 -565
rect -797 -605 -739 -599
rect -605 -565 -547 -559
rect -605 -599 -593 -565
rect -559 -599 -547 -565
rect -605 -605 -547 -599
rect -413 -565 -355 -559
rect -413 -599 -401 -565
rect -367 -599 -355 -565
rect -413 -605 -355 -599
rect -221 -565 -163 -559
rect -221 -599 -209 -565
rect -175 -599 -163 -565
rect -221 -605 -163 -599
rect -29 -565 29 -559
rect -29 -599 -17 -565
rect 17 -599 29 -565
rect -29 -605 29 -599
rect 163 -565 221 -559
rect 163 -599 175 -565
rect 209 -599 221 -565
rect 163 -605 221 -599
rect 355 -565 413 -559
rect 355 -599 367 -565
rect 401 -599 413 -565
rect 355 -605 413 -599
rect 547 -565 605 -559
rect 547 -599 559 -565
rect 593 -599 605 -565
rect 547 -605 605 -599
rect 739 -565 797 -559
rect 739 -599 751 -565
rect 785 -599 797 -565
rect 739 -605 797 -599
rect 931 -565 989 -559
rect 931 -599 943 -565
rect 977 -599 989 -565
rect 931 -605 989 -599
rect 1123 -565 1181 -559
rect 1123 -599 1135 -565
rect 1169 -599 1181 -565
rect 1123 -605 1181 -599
rect 1315 -565 1373 -559
rect 1315 -599 1327 -565
rect 1361 -599 1373 -565
rect 1315 -605 1373 -599
rect 1507 -565 1565 -559
rect 1507 -599 1519 -565
rect 1553 -599 1565 -565
rect 1507 -605 1565 -599
rect 1699 -565 1757 -559
rect 1699 -599 1711 -565
rect 1745 -599 1757 -565
rect 1699 -605 1757 -599
rect 1891 -565 1949 -559
rect 1891 -599 1903 -565
rect 1937 -599 1949 -565
rect 1891 -605 1949 -599
rect 2083 -565 2141 -559
rect 2083 -599 2095 -565
rect 2129 -599 2141 -565
rect 2083 -605 2141 -599
<< properties >>
string FIXED_BBOX -2274 -684 2274 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 2 nf 45 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
