magic
tech sky130A
magscale 1 2
timestamp 1645802395
<< metal4 >>
rect -951 3059 951 3100
rect -951 -3059 695 3059
rect 931 -3059 951 3059
rect -951 -3100 951 -3059
<< via4 >>
rect 695 -3059 931 3059
<< mimcap2 >>
rect -851 2960 349 3000
rect -851 -2960 -811 2960
rect 309 -2960 349 2960
rect -851 -3000 349 -2960
<< mimcap2contact >>
rect -811 -2960 309 2960
<< metal5 >>
rect 653 3059 973 3101
rect -835 2960 333 2984
rect -835 -2960 -811 2960
rect 309 -2960 333 2960
rect -835 -2984 333 -2960
rect 653 -3059 695 3059
rect 931 -3059 973 3059
rect 653 -3101 973 -3059
<< properties >>
string FIXED_BBOX -951 -3100 449 3100
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 6 l 30 val 373.68 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
