magic
tech sky130A
magscale 1 2
timestamp 1645541123
<< pwell >>
rect -1457 -2137 1457 2137
<< nmos >>
rect -1261 1127 -1061 1927
rect -1003 1127 -803 1927
rect -745 1127 -545 1927
rect -487 1127 -287 1927
rect -229 1127 -29 1927
rect 29 1127 229 1927
rect 287 1127 487 1927
rect 545 1127 745 1927
rect 803 1127 1003 1927
rect 1061 1127 1261 1927
rect -1261 109 -1061 909
rect -1003 109 -803 909
rect -745 109 -545 909
rect -487 109 -287 909
rect -229 109 -29 909
rect 29 109 229 909
rect 287 109 487 909
rect 545 109 745 909
rect 803 109 1003 909
rect 1061 109 1261 909
rect -1261 -909 -1061 -109
rect -1003 -909 -803 -109
rect -745 -909 -545 -109
rect -487 -909 -287 -109
rect -229 -909 -29 -109
rect 29 -909 229 -109
rect 287 -909 487 -109
rect 545 -909 745 -109
rect 803 -909 1003 -109
rect 1061 -909 1261 -109
rect -1261 -1927 -1061 -1127
rect -1003 -1927 -803 -1127
rect -745 -1927 -545 -1127
rect -487 -1927 -287 -1127
rect -229 -1927 -29 -1127
rect 29 -1927 229 -1127
rect 287 -1927 487 -1127
rect 545 -1927 745 -1127
rect 803 -1927 1003 -1127
rect 1061 -1927 1261 -1127
<< ndiff >>
rect -1319 1915 -1261 1927
rect -1319 1139 -1307 1915
rect -1273 1139 -1261 1915
rect -1319 1127 -1261 1139
rect -1061 1915 -1003 1927
rect -1061 1139 -1049 1915
rect -1015 1139 -1003 1915
rect -1061 1127 -1003 1139
rect -803 1915 -745 1927
rect -803 1139 -791 1915
rect -757 1139 -745 1915
rect -803 1127 -745 1139
rect -545 1915 -487 1927
rect -545 1139 -533 1915
rect -499 1139 -487 1915
rect -545 1127 -487 1139
rect -287 1915 -229 1927
rect -287 1139 -275 1915
rect -241 1139 -229 1915
rect -287 1127 -229 1139
rect -29 1915 29 1927
rect -29 1139 -17 1915
rect 17 1139 29 1915
rect -29 1127 29 1139
rect 229 1915 287 1927
rect 229 1139 241 1915
rect 275 1139 287 1915
rect 229 1127 287 1139
rect 487 1915 545 1927
rect 487 1139 499 1915
rect 533 1139 545 1915
rect 487 1127 545 1139
rect 745 1915 803 1927
rect 745 1139 757 1915
rect 791 1139 803 1915
rect 745 1127 803 1139
rect 1003 1915 1061 1927
rect 1003 1139 1015 1915
rect 1049 1139 1061 1915
rect 1003 1127 1061 1139
rect 1261 1915 1319 1927
rect 1261 1139 1273 1915
rect 1307 1139 1319 1915
rect 1261 1127 1319 1139
rect -1319 897 -1261 909
rect -1319 121 -1307 897
rect -1273 121 -1261 897
rect -1319 109 -1261 121
rect -1061 897 -1003 909
rect -1061 121 -1049 897
rect -1015 121 -1003 897
rect -1061 109 -1003 121
rect -803 897 -745 909
rect -803 121 -791 897
rect -757 121 -745 897
rect -803 109 -745 121
rect -545 897 -487 909
rect -545 121 -533 897
rect -499 121 -487 897
rect -545 109 -487 121
rect -287 897 -229 909
rect -287 121 -275 897
rect -241 121 -229 897
rect -287 109 -229 121
rect -29 897 29 909
rect -29 121 -17 897
rect 17 121 29 897
rect -29 109 29 121
rect 229 897 287 909
rect 229 121 241 897
rect 275 121 287 897
rect 229 109 287 121
rect 487 897 545 909
rect 487 121 499 897
rect 533 121 545 897
rect 487 109 545 121
rect 745 897 803 909
rect 745 121 757 897
rect 791 121 803 897
rect 745 109 803 121
rect 1003 897 1061 909
rect 1003 121 1015 897
rect 1049 121 1061 897
rect 1003 109 1061 121
rect 1261 897 1319 909
rect 1261 121 1273 897
rect 1307 121 1319 897
rect 1261 109 1319 121
rect -1319 -121 -1261 -109
rect -1319 -897 -1307 -121
rect -1273 -897 -1261 -121
rect -1319 -909 -1261 -897
rect -1061 -121 -1003 -109
rect -1061 -897 -1049 -121
rect -1015 -897 -1003 -121
rect -1061 -909 -1003 -897
rect -803 -121 -745 -109
rect -803 -897 -791 -121
rect -757 -897 -745 -121
rect -803 -909 -745 -897
rect -545 -121 -487 -109
rect -545 -897 -533 -121
rect -499 -897 -487 -121
rect -545 -909 -487 -897
rect -287 -121 -229 -109
rect -287 -897 -275 -121
rect -241 -897 -229 -121
rect -287 -909 -229 -897
rect -29 -121 29 -109
rect -29 -897 -17 -121
rect 17 -897 29 -121
rect -29 -909 29 -897
rect 229 -121 287 -109
rect 229 -897 241 -121
rect 275 -897 287 -121
rect 229 -909 287 -897
rect 487 -121 545 -109
rect 487 -897 499 -121
rect 533 -897 545 -121
rect 487 -909 545 -897
rect 745 -121 803 -109
rect 745 -897 757 -121
rect 791 -897 803 -121
rect 745 -909 803 -897
rect 1003 -121 1061 -109
rect 1003 -897 1015 -121
rect 1049 -897 1061 -121
rect 1003 -909 1061 -897
rect 1261 -121 1319 -109
rect 1261 -897 1273 -121
rect 1307 -897 1319 -121
rect 1261 -909 1319 -897
rect -1319 -1139 -1261 -1127
rect -1319 -1915 -1307 -1139
rect -1273 -1915 -1261 -1139
rect -1319 -1927 -1261 -1915
rect -1061 -1139 -1003 -1127
rect -1061 -1915 -1049 -1139
rect -1015 -1915 -1003 -1139
rect -1061 -1927 -1003 -1915
rect -803 -1139 -745 -1127
rect -803 -1915 -791 -1139
rect -757 -1915 -745 -1139
rect -803 -1927 -745 -1915
rect -545 -1139 -487 -1127
rect -545 -1915 -533 -1139
rect -499 -1915 -487 -1139
rect -545 -1927 -487 -1915
rect -287 -1139 -229 -1127
rect -287 -1915 -275 -1139
rect -241 -1915 -229 -1139
rect -287 -1927 -229 -1915
rect -29 -1139 29 -1127
rect -29 -1915 -17 -1139
rect 17 -1915 29 -1139
rect -29 -1927 29 -1915
rect 229 -1139 287 -1127
rect 229 -1915 241 -1139
rect 275 -1915 287 -1139
rect 229 -1927 287 -1915
rect 487 -1139 545 -1127
rect 487 -1915 499 -1139
rect 533 -1915 545 -1139
rect 487 -1927 545 -1915
rect 745 -1139 803 -1127
rect 745 -1915 757 -1139
rect 791 -1915 803 -1139
rect 745 -1927 803 -1915
rect 1003 -1139 1061 -1127
rect 1003 -1915 1015 -1139
rect 1049 -1915 1061 -1139
rect 1003 -1927 1061 -1915
rect 1261 -1139 1319 -1127
rect 1261 -1915 1273 -1139
rect 1307 -1915 1319 -1139
rect 1261 -1927 1319 -1915
<< ndiffc >>
rect -1307 1139 -1273 1915
rect -1049 1139 -1015 1915
rect -791 1139 -757 1915
rect -533 1139 -499 1915
rect -275 1139 -241 1915
rect -17 1139 17 1915
rect 241 1139 275 1915
rect 499 1139 533 1915
rect 757 1139 791 1915
rect 1015 1139 1049 1915
rect 1273 1139 1307 1915
rect -1307 121 -1273 897
rect -1049 121 -1015 897
rect -791 121 -757 897
rect -533 121 -499 897
rect -275 121 -241 897
rect -17 121 17 897
rect 241 121 275 897
rect 499 121 533 897
rect 757 121 791 897
rect 1015 121 1049 897
rect 1273 121 1307 897
rect -1307 -897 -1273 -121
rect -1049 -897 -1015 -121
rect -791 -897 -757 -121
rect -533 -897 -499 -121
rect -275 -897 -241 -121
rect -17 -897 17 -121
rect 241 -897 275 -121
rect 499 -897 533 -121
rect 757 -897 791 -121
rect 1015 -897 1049 -121
rect 1273 -897 1307 -121
rect -1307 -1915 -1273 -1139
rect -1049 -1915 -1015 -1139
rect -791 -1915 -757 -1139
rect -533 -1915 -499 -1139
rect -275 -1915 -241 -1139
rect -17 -1915 17 -1139
rect 241 -1915 275 -1139
rect 499 -1915 533 -1139
rect 757 -1915 791 -1139
rect 1015 -1915 1049 -1139
rect 1273 -1915 1307 -1139
<< psubdiff >>
rect -1421 2067 -1325 2101
rect 1325 2067 1421 2101
rect -1421 2005 -1387 2067
rect 1387 2005 1421 2067
rect -1421 -2067 -1387 -2005
rect 1387 -2067 1421 -2005
rect -1421 -2101 -1325 -2067
rect 1325 -2101 1421 -2067
<< psubdiffcont >>
rect -1325 2067 1325 2101
rect -1421 -2005 -1387 2005
rect 1387 -2005 1421 2005
rect -1325 -2101 1325 -2067
<< poly >>
rect -1261 1999 -1061 2015
rect -1261 1965 -1245 1999
rect -1077 1965 -1061 1999
rect -1261 1927 -1061 1965
rect -1003 1999 -803 2015
rect -1003 1965 -987 1999
rect -819 1965 -803 1999
rect -1003 1927 -803 1965
rect -745 1999 -545 2015
rect -745 1965 -729 1999
rect -561 1965 -545 1999
rect -745 1927 -545 1965
rect -487 1999 -287 2015
rect -487 1965 -471 1999
rect -303 1965 -287 1999
rect -487 1927 -287 1965
rect -229 1999 -29 2015
rect -229 1965 -213 1999
rect -45 1965 -29 1999
rect -229 1927 -29 1965
rect 29 1999 229 2015
rect 29 1965 45 1999
rect 213 1965 229 1999
rect 29 1927 229 1965
rect 287 1999 487 2015
rect 287 1965 303 1999
rect 471 1965 487 1999
rect 287 1927 487 1965
rect 545 1999 745 2015
rect 545 1965 561 1999
rect 729 1965 745 1999
rect 545 1927 745 1965
rect 803 1999 1003 2015
rect 803 1965 819 1999
rect 987 1965 1003 1999
rect 803 1927 1003 1965
rect 1061 1999 1261 2015
rect 1061 1965 1077 1999
rect 1245 1965 1261 1999
rect 1061 1927 1261 1965
rect -1261 1089 -1061 1127
rect -1261 1055 -1245 1089
rect -1077 1055 -1061 1089
rect -1261 1039 -1061 1055
rect -1003 1089 -803 1127
rect -1003 1055 -987 1089
rect -819 1055 -803 1089
rect -1003 1039 -803 1055
rect -745 1089 -545 1127
rect -745 1055 -729 1089
rect -561 1055 -545 1089
rect -745 1039 -545 1055
rect -487 1089 -287 1127
rect -487 1055 -471 1089
rect -303 1055 -287 1089
rect -487 1039 -287 1055
rect -229 1089 -29 1127
rect -229 1055 -213 1089
rect -45 1055 -29 1089
rect -229 1039 -29 1055
rect 29 1089 229 1127
rect 29 1055 45 1089
rect 213 1055 229 1089
rect 29 1039 229 1055
rect 287 1089 487 1127
rect 287 1055 303 1089
rect 471 1055 487 1089
rect 287 1039 487 1055
rect 545 1089 745 1127
rect 545 1055 561 1089
rect 729 1055 745 1089
rect 545 1039 745 1055
rect 803 1089 1003 1127
rect 803 1055 819 1089
rect 987 1055 1003 1089
rect 803 1039 1003 1055
rect 1061 1089 1261 1127
rect 1061 1055 1077 1089
rect 1245 1055 1261 1089
rect 1061 1039 1261 1055
rect -1261 981 -1061 997
rect -1261 947 -1245 981
rect -1077 947 -1061 981
rect -1261 909 -1061 947
rect -1003 981 -803 997
rect -1003 947 -987 981
rect -819 947 -803 981
rect -1003 909 -803 947
rect -745 981 -545 997
rect -745 947 -729 981
rect -561 947 -545 981
rect -745 909 -545 947
rect -487 981 -287 997
rect -487 947 -471 981
rect -303 947 -287 981
rect -487 909 -287 947
rect -229 981 -29 997
rect -229 947 -213 981
rect -45 947 -29 981
rect -229 909 -29 947
rect 29 981 229 997
rect 29 947 45 981
rect 213 947 229 981
rect 29 909 229 947
rect 287 981 487 997
rect 287 947 303 981
rect 471 947 487 981
rect 287 909 487 947
rect 545 981 745 997
rect 545 947 561 981
rect 729 947 745 981
rect 545 909 745 947
rect 803 981 1003 997
rect 803 947 819 981
rect 987 947 1003 981
rect 803 909 1003 947
rect 1061 981 1261 997
rect 1061 947 1077 981
rect 1245 947 1261 981
rect 1061 909 1261 947
rect -1261 71 -1061 109
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 109
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 109
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 109
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 109
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 109
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -109 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -109 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -109 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -109 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -109 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -109 1261 -71
rect -1261 -947 -1061 -909
rect -1261 -981 -1245 -947
rect -1077 -981 -1061 -947
rect -1261 -997 -1061 -981
rect -1003 -947 -803 -909
rect -1003 -981 -987 -947
rect -819 -981 -803 -947
rect -1003 -997 -803 -981
rect -745 -947 -545 -909
rect -745 -981 -729 -947
rect -561 -981 -545 -947
rect -745 -997 -545 -981
rect -487 -947 -287 -909
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -487 -997 -287 -981
rect -229 -947 -29 -909
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect -229 -997 -29 -981
rect 29 -947 229 -909
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 29 -997 229 -981
rect 287 -947 487 -909
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 287 -997 487 -981
rect 545 -947 745 -909
rect 545 -981 561 -947
rect 729 -981 745 -947
rect 545 -997 745 -981
rect 803 -947 1003 -909
rect 803 -981 819 -947
rect 987 -981 1003 -947
rect 803 -997 1003 -981
rect 1061 -947 1261 -909
rect 1061 -981 1077 -947
rect 1245 -981 1261 -947
rect 1061 -997 1261 -981
rect -1261 -1055 -1061 -1039
rect -1261 -1089 -1245 -1055
rect -1077 -1089 -1061 -1055
rect -1261 -1127 -1061 -1089
rect -1003 -1055 -803 -1039
rect -1003 -1089 -987 -1055
rect -819 -1089 -803 -1055
rect -1003 -1127 -803 -1089
rect -745 -1055 -545 -1039
rect -745 -1089 -729 -1055
rect -561 -1089 -545 -1055
rect -745 -1127 -545 -1089
rect -487 -1055 -287 -1039
rect -487 -1089 -471 -1055
rect -303 -1089 -287 -1055
rect -487 -1127 -287 -1089
rect -229 -1055 -29 -1039
rect -229 -1089 -213 -1055
rect -45 -1089 -29 -1055
rect -229 -1127 -29 -1089
rect 29 -1055 229 -1039
rect 29 -1089 45 -1055
rect 213 -1089 229 -1055
rect 29 -1127 229 -1089
rect 287 -1055 487 -1039
rect 287 -1089 303 -1055
rect 471 -1089 487 -1055
rect 287 -1127 487 -1089
rect 545 -1055 745 -1039
rect 545 -1089 561 -1055
rect 729 -1089 745 -1055
rect 545 -1127 745 -1089
rect 803 -1055 1003 -1039
rect 803 -1089 819 -1055
rect 987 -1089 1003 -1055
rect 803 -1127 1003 -1089
rect 1061 -1055 1261 -1039
rect 1061 -1089 1077 -1055
rect 1245 -1089 1261 -1055
rect 1061 -1127 1261 -1089
rect -1261 -1965 -1061 -1927
rect -1261 -1999 -1245 -1965
rect -1077 -1999 -1061 -1965
rect -1261 -2015 -1061 -1999
rect -1003 -1965 -803 -1927
rect -1003 -1999 -987 -1965
rect -819 -1999 -803 -1965
rect -1003 -2015 -803 -1999
rect -745 -1965 -545 -1927
rect -745 -1999 -729 -1965
rect -561 -1999 -545 -1965
rect -745 -2015 -545 -1999
rect -487 -1965 -287 -1927
rect -487 -1999 -471 -1965
rect -303 -1999 -287 -1965
rect -487 -2015 -287 -1999
rect -229 -1965 -29 -1927
rect -229 -1999 -213 -1965
rect -45 -1999 -29 -1965
rect -229 -2015 -29 -1999
rect 29 -1965 229 -1927
rect 29 -1999 45 -1965
rect 213 -1999 229 -1965
rect 29 -2015 229 -1999
rect 287 -1965 487 -1927
rect 287 -1999 303 -1965
rect 471 -1999 487 -1965
rect 287 -2015 487 -1999
rect 545 -1965 745 -1927
rect 545 -1999 561 -1965
rect 729 -1999 745 -1965
rect 545 -2015 745 -1999
rect 803 -1965 1003 -1927
rect 803 -1999 819 -1965
rect 987 -1999 1003 -1965
rect 803 -2015 1003 -1999
rect 1061 -1965 1261 -1927
rect 1061 -1999 1077 -1965
rect 1245 -1999 1261 -1965
rect 1061 -2015 1261 -1999
<< polycont >>
rect -1245 1965 -1077 1999
rect -987 1965 -819 1999
rect -729 1965 -561 1999
rect -471 1965 -303 1999
rect -213 1965 -45 1999
rect 45 1965 213 1999
rect 303 1965 471 1999
rect 561 1965 729 1999
rect 819 1965 987 1999
rect 1077 1965 1245 1999
rect -1245 1055 -1077 1089
rect -987 1055 -819 1089
rect -729 1055 -561 1089
rect -471 1055 -303 1089
rect -213 1055 -45 1089
rect 45 1055 213 1089
rect 303 1055 471 1089
rect 561 1055 729 1089
rect 819 1055 987 1089
rect 1077 1055 1245 1089
rect -1245 947 -1077 981
rect -987 947 -819 981
rect -729 947 -561 981
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect 561 947 729 981
rect 819 947 987 981
rect 1077 947 1245 981
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect -1245 -981 -1077 -947
rect -987 -981 -819 -947
rect -729 -981 -561 -947
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
rect 561 -981 729 -947
rect 819 -981 987 -947
rect 1077 -981 1245 -947
rect -1245 -1089 -1077 -1055
rect -987 -1089 -819 -1055
rect -729 -1089 -561 -1055
rect -471 -1089 -303 -1055
rect -213 -1089 -45 -1055
rect 45 -1089 213 -1055
rect 303 -1089 471 -1055
rect 561 -1089 729 -1055
rect 819 -1089 987 -1055
rect 1077 -1089 1245 -1055
rect -1245 -1999 -1077 -1965
rect -987 -1999 -819 -1965
rect -729 -1999 -561 -1965
rect -471 -1999 -303 -1965
rect -213 -1999 -45 -1965
rect 45 -1999 213 -1965
rect 303 -1999 471 -1965
rect 561 -1999 729 -1965
rect 819 -1999 987 -1965
rect 1077 -1999 1245 -1965
<< locali >>
rect -1421 2067 -1325 2101
rect 1325 2067 1421 2101
rect -1421 2005 -1387 2067
rect 1387 2005 1421 2067
rect -1261 1965 -1245 1999
rect -1077 1965 -1061 1999
rect -1003 1965 -987 1999
rect -819 1965 -803 1999
rect -745 1965 -729 1999
rect -561 1965 -545 1999
rect -487 1965 -471 1999
rect -303 1965 -287 1999
rect -229 1965 -213 1999
rect -45 1965 -29 1999
rect 29 1965 45 1999
rect 213 1965 229 1999
rect 287 1965 303 1999
rect 471 1965 487 1999
rect 545 1965 561 1999
rect 729 1965 745 1999
rect 803 1965 819 1999
rect 987 1965 1003 1999
rect 1061 1965 1077 1999
rect 1245 1965 1261 1999
rect -1307 1915 -1273 1931
rect -1307 1123 -1273 1139
rect -1049 1915 -1015 1931
rect -1049 1123 -1015 1139
rect -791 1915 -757 1931
rect -791 1123 -757 1139
rect -533 1915 -499 1931
rect -533 1123 -499 1139
rect -275 1915 -241 1931
rect -275 1123 -241 1139
rect -17 1915 17 1931
rect -17 1123 17 1139
rect 241 1915 275 1931
rect 241 1123 275 1139
rect 499 1915 533 1931
rect 499 1123 533 1139
rect 757 1915 791 1931
rect 757 1123 791 1139
rect 1015 1915 1049 1931
rect 1015 1123 1049 1139
rect 1273 1915 1307 1931
rect 1273 1123 1307 1139
rect -1261 1055 -1245 1089
rect -1077 1055 -1061 1089
rect -1003 1055 -987 1089
rect -819 1055 -803 1089
rect -745 1055 -729 1089
rect -561 1055 -545 1089
rect -487 1055 -471 1089
rect -303 1055 -287 1089
rect -229 1055 -213 1089
rect -45 1055 -29 1089
rect 29 1055 45 1089
rect 213 1055 229 1089
rect 287 1055 303 1089
rect 471 1055 487 1089
rect 545 1055 561 1089
rect 729 1055 745 1089
rect 803 1055 819 1089
rect 987 1055 1003 1089
rect 1061 1055 1077 1089
rect 1245 1055 1261 1089
rect -1261 947 -1245 981
rect -1077 947 -1061 981
rect -1003 947 -987 981
rect -819 947 -803 981
rect -745 947 -729 981
rect -561 947 -545 981
rect -487 947 -471 981
rect -303 947 -287 981
rect -229 947 -213 981
rect -45 947 -29 981
rect 29 947 45 981
rect 213 947 229 981
rect 287 947 303 981
rect 471 947 487 981
rect 545 947 561 981
rect 729 947 745 981
rect 803 947 819 981
rect 987 947 1003 981
rect 1061 947 1077 981
rect 1245 947 1261 981
rect -1307 897 -1273 913
rect -1307 105 -1273 121
rect -1049 897 -1015 913
rect -1049 105 -1015 121
rect -791 897 -757 913
rect -791 105 -757 121
rect -533 897 -499 913
rect -533 105 -499 121
rect -275 897 -241 913
rect -275 105 -241 121
rect -17 897 17 913
rect -17 105 17 121
rect 241 897 275 913
rect 241 105 275 121
rect 499 897 533 913
rect 499 105 533 121
rect 757 897 791 913
rect 757 105 791 121
rect 1015 897 1049 913
rect 1015 105 1049 121
rect 1273 897 1307 913
rect 1273 105 1307 121
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect -1307 -121 -1273 -105
rect -1307 -913 -1273 -897
rect -1049 -121 -1015 -105
rect -1049 -913 -1015 -897
rect -791 -121 -757 -105
rect -791 -913 -757 -897
rect -533 -121 -499 -105
rect -533 -913 -499 -897
rect -275 -121 -241 -105
rect -275 -913 -241 -897
rect -17 -121 17 -105
rect -17 -913 17 -897
rect 241 -121 275 -105
rect 241 -913 275 -897
rect 499 -121 533 -105
rect 499 -913 533 -897
rect 757 -121 791 -105
rect 757 -913 791 -897
rect 1015 -121 1049 -105
rect 1015 -913 1049 -897
rect 1273 -121 1307 -105
rect 1273 -913 1307 -897
rect -1261 -981 -1245 -947
rect -1077 -981 -1061 -947
rect -1003 -981 -987 -947
rect -819 -981 -803 -947
rect -745 -981 -729 -947
rect -561 -981 -545 -947
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 545 -981 561 -947
rect 729 -981 745 -947
rect 803 -981 819 -947
rect 987 -981 1003 -947
rect 1061 -981 1077 -947
rect 1245 -981 1261 -947
rect -1261 -1089 -1245 -1055
rect -1077 -1089 -1061 -1055
rect -1003 -1089 -987 -1055
rect -819 -1089 -803 -1055
rect -745 -1089 -729 -1055
rect -561 -1089 -545 -1055
rect -487 -1089 -471 -1055
rect -303 -1089 -287 -1055
rect -229 -1089 -213 -1055
rect -45 -1089 -29 -1055
rect 29 -1089 45 -1055
rect 213 -1089 229 -1055
rect 287 -1089 303 -1055
rect 471 -1089 487 -1055
rect 545 -1089 561 -1055
rect 729 -1089 745 -1055
rect 803 -1089 819 -1055
rect 987 -1089 1003 -1055
rect 1061 -1089 1077 -1055
rect 1245 -1089 1261 -1055
rect -1307 -1139 -1273 -1123
rect -1307 -1931 -1273 -1915
rect -1049 -1139 -1015 -1123
rect -1049 -1931 -1015 -1915
rect -791 -1139 -757 -1123
rect -791 -1931 -757 -1915
rect -533 -1139 -499 -1123
rect -533 -1931 -499 -1915
rect -275 -1139 -241 -1123
rect -275 -1931 -241 -1915
rect -17 -1139 17 -1123
rect -17 -1931 17 -1915
rect 241 -1139 275 -1123
rect 241 -1931 275 -1915
rect 499 -1139 533 -1123
rect 499 -1931 533 -1915
rect 757 -1139 791 -1123
rect 757 -1931 791 -1915
rect 1015 -1139 1049 -1123
rect 1015 -1931 1049 -1915
rect 1273 -1139 1307 -1123
rect 1273 -1931 1307 -1915
rect -1261 -1999 -1245 -1965
rect -1077 -1999 -1061 -1965
rect -1003 -1999 -987 -1965
rect -819 -1999 -803 -1965
rect -745 -1999 -729 -1965
rect -561 -1999 -545 -1965
rect -487 -1999 -471 -1965
rect -303 -1999 -287 -1965
rect -229 -1999 -213 -1965
rect -45 -1999 -29 -1965
rect 29 -1999 45 -1965
rect 213 -1999 229 -1965
rect 287 -1999 303 -1965
rect 471 -1999 487 -1965
rect 545 -1999 561 -1965
rect 729 -1999 745 -1965
rect 803 -1999 819 -1965
rect 987 -1999 1003 -1965
rect 1061 -1999 1077 -1965
rect 1245 -1999 1261 -1965
rect -1421 -2067 -1387 -2005
rect 1387 -2067 1421 -2005
rect -1421 -2101 -1325 -2067
rect 1325 -2101 1421 -2067
<< viali >>
rect -1245 1965 -1077 1999
rect -987 1965 -819 1999
rect -729 1965 -561 1999
rect -471 1965 -303 1999
rect -213 1965 -45 1999
rect 45 1965 213 1999
rect 303 1965 471 1999
rect 561 1965 729 1999
rect 819 1965 987 1999
rect 1077 1965 1245 1999
rect -1307 1139 -1273 1915
rect -1049 1139 -1015 1915
rect -791 1139 -757 1915
rect -533 1139 -499 1915
rect -275 1139 -241 1915
rect -17 1139 17 1915
rect 241 1139 275 1915
rect 499 1139 533 1915
rect 757 1139 791 1915
rect 1015 1139 1049 1915
rect 1273 1139 1307 1915
rect -1245 1055 -1077 1089
rect -987 1055 -819 1089
rect -729 1055 -561 1089
rect -471 1055 -303 1089
rect -213 1055 -45 1089
rect 45 1055 213 1089
rect 303 1055 471 1089
rect 561 1055 729 1089
rect 819 1055 987 1089
rect 1077 1055 1245 1089
rect -1245 947 -1077 981
rect -987 947 -819 981
rect -729 947 -561 981
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect 561 947 729 981
rect 819 947 987 981
rect 1077 947 1245 981
rect -1307 121 -1273 897
rect -1049 121 -1015 897
rect -791 121 -757 897
rect -533 121 -499 897
rect -275 121 -241 897
rect -17 121 17 897
rect 241 121 275 897
rect 499 121 533 897
rect 757 121 791 897
rect 1015 121 1049 897
rect 1273 121 1307 897
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect -1307 -897 -1273 -121
rect -1049 -897 -1015 -121
rect -791 -897 -757 -121
rect -533 -897 -499 -121
rect -275 -897 -241 -121
rect -17 -897 17 -121
rect 241 -897 275 -121
rect 499 -897 533 -121
rect 757 -897 791 -121
rect 1015 -897 1049 -121
rect 1273 -897 1307 -121
rect -1245 -981 -1077 -947
rect -987 -981 -819 -947
rect -729 -981 -561 -947
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
rect 561 -981 729 -947
rect 819 -981 987 -947
rect 1077 -981 1245 -947
rect -1245 -1089 -1077 -1055
rect -987 -1089 -819 -1055
rect -729 -1089 -561 -1055
rect -471 -1089 -303 -1055
rect -213 -1089 -45 -1055
rect 45 -1089 213 -1055
rect 303 -1089 471 -1055
rect 561 -1089 729 -1055
rect 819 -1089 987 -1055
rect 1077 -1089 1245 -1055
rect -1307 -1915 -1273 -1139
rect -1049 -1915 -1015 -1139
rect -791 -1915 -757 -1139
rect -533 -1915 -499 -1139
rect -275 -1915 -241 -1139
rect -17 -1915 17 -1139
rect 241 -1915 275 -1139
rect 499 -1915 533 -1139
rect 757 -1915 791 -1139
rect 1015 -1915 1049 -1139
rect 1273 -1915 1307 -1139
rect -1245 -1999 -1077 -1965
rect -987 -1999 -819 -1965
rect -729 -1999 -561 -1965
rect -471 -1999 -303 -1965
rect -213 -1999 -45 -1965
rect 45 -1999 213 -1965
rect 303 -1999 471 -1965
rect 561 -1999 729 -1965
rect 819 -1999 987 -1965
rect 1077 -1999 1245 -1965
<< metal1 >>
rect -1257 1999 -1065 2005
rect -1257 1965 -1245 1999
rect -1077 1965 -1065 1999
rect -1257 1959 -1065 1965
rect -999 1999 -807 2005
rect -999 1965 -987 1999
rect -819 1965 -807 1999
rect -999 1959 -807 1965
rect -741 1999 -549 2005
rect -741 1965 -729 1999
rect -561 1965 -549 1999
rect -741 1959 -549 1965
rect -483 1999 -291 2005
rect -483 1965 -471 1999
rect -303 1965 -291 1999
rect -483 1959 -291 1965
rect -225 1999 -33 2005
rect -225 1965 -213 1999
rect -45 1965 -33 1999
rect -225 1959 -33 1965
rect 33 1999 225 2005
rect 33 1965 45 1999
rect 213 1965 225 1999
rect 33 1959 225 1965
rect 291 1999 483 2005
rect 291 1965 303 1999
rect 471 1965 483 1999
rect 291 1959 483 1965
rect 549 1999 741 2005
rect 549 1965 561 1999
rect 729 1965 741 1999
rect 549 1959 741 1965
rect 807 1999 999 2005
rect 807 1965 819 1999
rect 987 1965 999 1999
rect 807 1959 999 1965
rect 1065 1999 1257 2005
rect 1065 1965 1077 1999
rect 1245 1965 1257 1999
rect 1065 1959 1257 1965
rect -1313 1915 -1267 1927
rect -1313 1139 -1307 1915
rect -1273 1139 -1267 1915
rect -1313 1127 -1267 1139
rect -1055 1915 -1009 1927
rect -1055 1139 -1049 1915
rect -1015 1139 -1009 1915
rect -1055 1127 -1009 1139
rect -797 1915 -751 1927
rect -797 1139 -791 1915
rect -757 1139 -751 1915
rect -797 1127 -751 1139
rect -539 1915 -493 1927
rect -539 1139 -533 1915
rect -499 1139 -493 1915
rect -539 1127 -493 1139
rect -281 1915 -235 1927
rect -281 1139 -275 1915
rect -241 1139 -235 1915
rect -281 1127 -235 1139
rect -23 1915 23 1927
rect -23 1139 -17 1915
rect 17 1139 23 1915
rect -23 1127 23 1139
rect 235 1915 281 1927
rect 235 1139 241 1915
rect 275 1139 281 1915
rect 235 1127 281 1139
rect 493 1915 539 1927
rect 493 1139 499 1915
rect 533 1139 539 1915
rect 493 1127 539 1139
rect 751 1915 797 1927
rect 751 1139 757 1915
rect 791 1139 797 1915
rect 751 1127 797 1139
rect 1009 1915 1055 1927
rect 1009 1139 1015 1915
rect 1049 1139 1055 1915
rect 1009 1127 1055 1139
rect 1267 1915 1313 1927
rect 1267 1139 1273 1915
rect 1307 1139 1313 1915
rect 1267 1127 1313 1139
rect -1257 1089 -1065 1095
rect -1257 1055 -1245 1089
rect -1077 1055 -1065 1089
rect -1257 1049 -1065 1055
rect -999 1089 -807 1095
rect -999 1055 -987 1089
rect -819 1055 -807 1089
rect -999 1049 -807 1055
rect -741 1089 -549 1095
rect -741 1055 -729 1089
rect -561 1055 -549 1089
rect -741 1049 -549 1055
rect -483 1089 -291 1095
rect -483 1055 -471 1089
rect -303 1055 -291 1089
rect -483 1049 -291 1055
rect -225 1089 -33 1095
rect -225 1055 -213 1089
rect -45 1055 -33 1089
rect -225 1049 -33 1055
rect 33 1089 225 1095
rect 33 1055 45 1089
rect 213 1055 225 1089
rect 33 1049 225 1055
rect 291 1089 483 1095
rect 291 1055 303 1089
rect 471 1055 483 1089
rect 291 1049 483 1055
rect 549 1089 741 1095
rect 549 1055 561 1089
rect 729 1055 741 1089
rect 549 1049 741 1055
rect 807 1089 999 1095
rect 807 1055 819 1089
rect 987 1055 999 1089
rect 807 1049 999 1055
rect 1065 1089 1257 1095
rect 1065 1055 1077 1089
rect 1245 1055 1257 1089
rect 1065 1049 1257 1055
rect -1257 981 -1065 987
rect -1257 947 -1245 981
rect -1077 947 -1065 981
rect -1257 941 -1065 947
rect -999 981 -807 987
rect -999 947 -987 981
rect -819 947 -807 981
rect -999 941 -807 947
rect -741 981 -549 987
rect -741 947 -729 981
rect -561 947 -549 981
rect -741 941 -549 947
rect -483 981 -291 987
rect -483 947 -471 981
rect -303 947 -291 981
rect -483 941 -291 947
rect -225 981 -33 987
rect -225 947 -213 981
rect -45 947 -33 981
rect -225 941 -33 947
rect 33 981 225 987
rect 33 947 45 981
rect 213 947 225 981
rect 33 941 225 947
rect 291 981 483 987
rect 291 947 303 981
rect 471 947 483 981
rect 291 941 483 947
rect 549 981 741 987
rect 549 947 561 981
rect 729 947 741 981
rect 549 941 741 947
rect 807 981 999 987
rect 807 947 819 981
rect 987 947 999 981
rect 807 941 999 947
rect 1065 981 1257 987
rect 1065 947 1077 981
rect 1245 947 1257 981
rect 1065 941 1257 947
rect -1313 897 -1267 909
rect -1313 121 -1307 897
rect -1273 121 -1267 897
rect -1313 109 -1267 121
rect -1055 897 -1009 909
rect -1055 121 -1049 897
rect -1015 121 -1009 897
rect -1055 109 -1009 121
rect -797 897 -751 909
rect -797 121 -791 897
rect -757 121 -751 897
rect -797 109 -751 121
rect -539 897 -493 909
rect -539 121 -533 897
rect -499 121 -493 897
rect -539 109 -493 121
rect -281 897 -235 909
rect -281 121 -275 897
rect -241 121 -235 897
rect -281 109 -235 121
rect -23 897 23 909
rect -23 121 -17 897
rect 17 121 23 897
rect -23 109 23 121
rect 235 897 281 909
rect 235 121 241 897
rect 275 121 281 897
rect 235 109 281 121
rect 493 897 539 909
rect 493 121 499 897
rect 533 121 539 897
rect 493 109 539 121
rect 751 897 797 909
rect 751 121 757 897
rect 791 121 797 897
rect 751 109 797 121
rect 1009 897 1055 909
rect 1009 121 1015 897
rect 1049 121 1055 897
rect 1009 109 1055 121
rect 1267 897 1313 909
rect 1267 121 1273 897
rect 1307 121 1313 897
rect 1267 109 1313 121
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect -1313 -121 -1267 -109
rect -1313 -897 -1307 -121
rect -1273 -897 -1267 -121
rect -1313 -909 -1267 -897
rect -1055 -121 -1009 -109
rect -1055 -897 -1049 -121
rect -1015 -897 -1009 -121
rect -1055 -909 -1009 -897
rect -797 -121 -751 -109
rect -797 -897 -791 -121
rect -757 -897 -751 -121
rect -797 -909 -751 -897
rect -539 -121 -493 -109
rect -539 -897 -533 -121
rect -499 -897 -493 -121
rect -539 -909 -493 -897
rect -281 -121 -235 -109
rect -281 -897 -275 -121
rect -241 -897 -235 -121
rect -281 -909 -235 -897
rect -23 -121 23 -109
rect -23 -897 -17 -121
rect 17 -897 23 -121
rect -23 -909 23 -897
rect 235 -121 281 -109
rect 235 -897 241 -121
rect 275 -897 281 -121
rect 235 -909 281 -897
rect 493 -121 539 -109
rect 493 -897 499 -121
rect 533 -897 539 -121
rect 493 -909 539 -897
rect 751 -121 797 -109
rect 751 -897 757 -121
rect 791 -897 797 -121
rect 751 -909 797 -897
rect 1009 -121 1055 -109
rect 1009 -897 1015 -121
rect 1049 -897 1055 -121
rect 1009 -909 1055 -897
rect 1267 -121 1313 -109
rect 1267 -897 1273 -121
rect 1307 -897 1313 -121
rect 1267 -909 1313 -897
rect -1257 -947 -1065 -941
rect -1257 -981 -1245 -947
rect -1077 -981 -1065 -947
rect -1257 -987 -1065 -981
rect -999 -947 -807 -941
rect -999 -981 -987 -947
rect -819 -981 -807 -947
rect -999 -987 -807 -981
rect -741 -947 -549 -941
rect -741 -981 -729 -947
rect -561 -981 -549 -947
rect -741 -987 -549 -981
rect -483 -947 -291 -941
rect -483 -981 -471 -947
rect -303 -981 -291 -947
rect -483 -987 -291 -981
rect -225 -947 -33 -941
rect -225 -981 -213 -947
rect -45 -981 -33 -947
rect -225 -987 -33 -981
rect 33 -947 225 -941
rect 33 -981 45 -947
rect 213 -981 225 -947
rect 33 -987 225 -981
rect 291 -947 483 -941
rect 291 -981 303 -947
rect 471 -981 483 -947
rect 291 -987 483 -981
rect 549 -947 741 -941
rect 549 -981 561 -947
rect 729 -981 741 -947
rect 549 -987 741 -981
rect 807 -947 999 -941
rect 807 -981 819 -947
rect 987 -981 999 -947
rect 807 -987 999 -981
rect 1065 -947 1257 -941
rect 1065 -981 1077 -947
rect 1245 -981 1257 -947
rect 1065 -987 1257 -981
rect -1257 -1055 -1065 -1049
rect -1257 -1089 -1245 -1055
rect -1077 -1089 -1065 -1055
rect -1257 -1095 -1065 -1089
rect -999 -1055 -807 -1049
rect -999 -1089 -987 -1055
rect -819 -1089 -807 -1055
rect -999 -1095 -807 -1089
rect -741 -1055 -549 -1049
rect -741 -1089 -729 -1055
rect -561 -1089 -549 -1055
rect -741 -1095 -549 -1089
rect -483 -1055 -291 -1049
rect -483 -1089 -471 -1055
rect -303 -1089 -291 -1055
rect -483 -1095 -291 -1089
rect -225 -1055 -33 -1049
rect -225 -1089 -213 -1055
rect -45 -1089 -33 -1055
rect -225 -1095 -33 -1089
rect 33 -1055 225 -1049
rect 33 -1089 45 -1055
rect 213 -1089 225 -1055
rect 33 -1095 225 -1089
rect 291 -1055 483 -1049
rect 291 -1089 303 -1055
rect 471 -1089 483 -1055
rect 291 -1095 483 -1089
rect 549 -1055 741 -1049
rect 549 -1089 561 -1055
rect 729 -1089 741 -1055
rect 549 -1095 741 -1089
rect 807 -1055 999 -1049
rect 807 -1089 819 -1055
rect 987 -1089 999 -1055
rect 807 -1095 999 -1089
rect 1065 -1055 1257 -1049
rect 1065 -1089 1077 -1055
rect 1245 -1089 1257 -1055
rect 1065 -1095 1257 -1089
rect -1313 -1139 -1267 -1127
rect -1313 -1915 -1307 -1139
rect -1273 -1915 -1267 -1139
rect -1313 -1927 -1267 -1915
rect -1055 -1139 -1009 -1127
rect -1055 -1915 -1049 -1139
rect -1015 -1915 -1009 -1139
rect -1055 -1927 -1009 -1915
rect -797 -1139 -751 -1127
rect -797 -1915 -791 -1139
rect -757 -1915 -751 -1139
rect -797 -1927 -751 -1915
rect -539 -1139 -493 -1127
rect -539 -1915 -533 -1139
rect -499 -1915 -493 -1139
rect -539 -1927 -493 -1915
rect -281 -1139 -235 -1127
rect -281 -1915 -275 -1139
rect -241 -1915 -235 -1139
rect -281 -1927 -235 -1915
rect -23 -1139 23 -1127
rect -23 -1915 -17 -1139
rect 17 -1915 23 -1139
rect -23 -1927 23 -1915
rect 235 -1139 281 -1127
rect 235 -1915 241 -1139
rect 275 -1915 281 -1139
rect 235 -1927 281 -1915
rect 493 -1139 539 -1127
rect 493 -1915 499 -1139
rect 533 -1915 539 -1139
rect 493 -1927 539 -1915
rect 751 -1139 797 -1127
rect 751 -1915 757 -1139
rect 791 -1915 797 -1139
rect 751 -1927 797 -1915
rect 1009 -1139 1055 -1127
rect 1009 -1915 1015 -1139
rect 1049 -1915 1055 -1139
rect 1009 -1927 1055 -1915
rect 1267 -1139 1313 -1127
rect 1267 -1915 1273 -1139
rect 1307 -1915 1313 -1139
rect 1267 -1927 1313 -1915
rect -1257 -1965 -1065 -1959
rect -1257 -1999 -1245 -1965
rect -1077 -1999 -1065 -1965
rect -1257 -2005 -1065 -1999
rect -999 -1965 -807 -1959
rect -999 -1999 -987 -1965
rect -819 -1999 -807 -1965
rect -999 -2005 -807 -1999
rect -741 -1965 -549 -1959
rect -741 -1999 -729 -1965
rect -561 -1999 -549 -1965
rect -741 -2005 -549 -1999
rect -483 -1965 -291 -1959
rect -483 -1999 -471 -1965
rect -303 -1999 -291 -1965
rect -483 -2005 -291 -1999
rect -225 -1965 -33 -1959
rect -225 -1999 -213 -1965
rect -45 -1999 -33 -1965
rect -225 -2005 -33 -1999
rect 33 -1965 225 -1959
rect 33 -1999 45 -1965
rect 213 -1999 225 -1965
rect 33 -2005 225 -1999
rect 291 -1965 483 -1959
rect 291 -1999 303 -1965
rect 471 -1999 483 -1965
rect 291 -2005 483 -1999
rect 549 -1965 741 -1959
rect 549 -1999 561 -1965
rect 729 -1999 741 -1965
rect 549 -2005 741 -1999
rect 807 -1965 999 -1959
rect 807 -1999 819 -1965
rect 987 -1999 999 -1965
rect 807 -2005 999 -1999
rect 1065 -1965 1257 -1959
rect 1065 -1999 1077 -1965
rect 1245 -1999 1257 -1965
rect 1065 -2005 1257 -1999
<< properties >>
string FIXED_BBOX -1404 -2084 1404 2084
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 1 m 4 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
