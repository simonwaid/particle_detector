magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< error_p >>
rect -269 281 -211 287
rect -77 281 -19 287
rect 115 281 173 287
rect 307 281 365 287
rect -269 247 -257 281
rect -77 247 -65 281
rect 115 247 127 281
rect 307 247 319 281
rect -269 241 -211 247
rect -77 241 -19 247
rect 115 241 173 247
rect 307 241 365 247
rect -365 -247 -307 -241
rect -173 -247 -115 -241
rect 19 -247 77 -241
rect 211 -247 269 -241
rect -365 -281 -353 -247
rect -173 -281 -161 -247
rect 19 -281 31 -247
rect 211 -281 223 -247
rect -365 -287 -307 -281
rect -173 -287 -115 -281
rect 19 -287 77 -281
rect 211 -287 269 -281
<< nwell >>
rect -551 -419 551 419
<< pmos >>
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
<< pdiff >>
rect -413 188 -351 200
rect -413 -188 -401 188
rect -367 -188 -351 188
rect -413 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 413 200
rect 351 -188 367 188
rect 401 -188 413 188
rect 351 -200 413 -188
<< pdiffc >>
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
<< nsubdiff >>
rect -515 349 -419 383
rect 419 349 515 383
rect -515 287 -481 349
rect 481 287 515 349
rect -515 -349 -481 -287
rect 481 -349 515 -287
rect -515 -383 -419 -349
rect 419 -383 515 -349
<< nsubdiffcont >>
rect -419 349 419 383
rect -515 -287 -481 287
rect 481 -287 515 287
rect -419 -383 419 -349
<< poly >>
rect -273 281 -207 297
rect -273 247 -257 281
rect -223 247 -207 281
rect -273 231 -207 247
rect -81 281 -15 297
rect -81 247 -65 281
rect -31 247 -15 281
rect -81 231 -15 247
rect 111 281 177 297
rect 111 247 127 281
rect 161 247 177 281
rect 111 231 177 247
rect 303 281 369 297
rect 303 247 319 281
rect 353 247 369 281
rect 303 231 369 247
rect -351 200 -321 226
rect -255 200 -225 231
rect -159 200 -129 226
rect -63 200 -33 231
rect 33 200 63 226
rect 129 200 159 231
rect 225 200 255 226
rect 321 200 351 231
rect -351 -231 -321 -200
rect -255 -226 -225 -200
rect -159 -231 -129 -200
rect -63 -226 -33 -200
rect 33 -231 63 -200
rect 129 -226 159 -200
rect 225 -231 255 -200
rect 321 -226 351 -200
rect -369 -247 -303 -231
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -369 -297 -303 -281
rect -177 -247 -111 -231
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect -177 -297 -111 -281
rect 15 -247 81 -231
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 15 -297 81 -281
rect 207 -247 273 -231
rect 207 -281 223 -247
rect 257 -281 273 -247
rect 207 -297 273 -281
<< polycont >>
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
<< locali >>
rect -515 349 -419 383
rect 419 349 515 383
rect -515 287 -481 349
rect 481 287 515 349
rect -273 247 -257 281
rect -223 247 -207 281
rect -81 247 -65 281
rect -31 247 -15 281
rect 111 247 127 281
rect 161 247 177 281
rect 303 247 319 281
rect 353 247 369 281
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 207 -281 223 -247
rect 257 -281 273 -247
rect -515 -349 -481 -287
rect 481 -349 515 -287
rect -515 -383 -419 -349
rect 419 -383 515 -349
<< viali >>
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
<< metal1 >>
rect -269 281 -211 287
rect -269 247 -257 281
rect -223 247 -211 281
rect -269 241 -211 247
rect -77 281 -19 287
rect -77 247 -65 281
rect -31 247 -19 281
rect -77 241 -19 247
rect 115 281 173 287
rect 115 247 127 281
rect 161 247 173 281
rect 115 241 173 247
rect 307 281 365 287
rect 307 247 319 281
rect 353 247 365 281
rect 307 241 365 247
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect -365 -247 -307 -241
rect -365 -281 -353 -247
rect -319 -281 -307 -247
rect -365 -287 -307 -281
rect -173 -247 -115 -241
rect -173 -281 -161 -247
rect -127 -281 -115 -247
rect -173 -287 -115 -281
rect 19 -247 77 -241
rect 19 -281 31 -247
rect 65 -281 77 -247
rect 19 -287 77 -281
rect 211 -247 269 -241
rect 211 -281 223 -247
rect 257 -281 269 -247
rect 211 -287 269 -281
<< properties >>
string FIXED_BBOX -498 -366 498 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
