magic
tech sky130A
magscale 1 2
timestamp 1654756835
<< nwell >>
rect -6340 4280 -6170 4450
rect -1290 4230 -1060 4450
rect 8150 4270 8320 4450
<< pwell >>
rect 4450 1180 4770 1210
rect 4960 1180 7980 1210
rect 4460 670 4780 700
rect 4960 670 7970 700
<< locali >>
rect 1420 1400 1520 2140
rect 850 1310 2090 1400
rect 1430 560 1510 1310
rect -640 -960 -530 -890
rect -630 -1600 -510 -1530
rect -110 -1590 -30 -1520
<< viali >>
rect 1360 4400 1660 4510
rect 6420 2590 6990 2690
rect -5630 -1530 -5550 -1370
rect -30 -1670 40 -1490
<< metal1 >>
rect -4170 6580 -3860 6630
rect -2820 6580 -2510 6630
rect 5210 6580 5610 6630
rect 6540 6580 6940 6630
rect 10120 6580 10450 6630
rect 11200 6580 11530 6630
rect -5000 5770 -4950 6070
rect -4140 6050 -3830 6100
rect -3660 5770 -3610 6070
rect -2790 6050 -2480 6100
rect -2320 5790 -2270 6090
rect 4140 6050 7980 6100
rect 4380 5730 4430 6050
rect 5720 5730 5770 6050
rect 7060 5730 7110 6050
rect 9810 5770 9870 6070
rect 10130 6050 10460 6100
rect 10900 5780 10960 6080
rect 11230 6050 11560 6100
rect 11990 5780 12050 6080
rect -4150 4940 -3860 4990
rect -2790 4940 -2500 4990
rect 5210 4940 5610 4990
rect 6550 4940 6950 4990
rect 10120 4940 10450 4990
rect 11230 4940 11560 4990
rect 830 4590 840 4750
rect 1440 4590 1450 4750
rect 1820 4580 1830 4750
rect 2310 4580 2320 4750
rect 1348 4510 1672 4516
rect -5000 4150 -4950 4450
rect -4160 4410 -3870 4460
rect -3660 4140 -3610 4440
rect -2810 4410 -2520 4460
rect -2320 4140 -2270 4440
rect 1348 4394 1360 4510
rect 1350 4340 1360 4394
rect 1660 4394 1672 4510
rect 4140 4410 7980 4460
rect 1660 4340 1670 4394
rect 4380 4090 4430 4410
rect 5720 4090 5770 4410
rect 7060 4090 7110 4410
rect 9810 4150 9870 4450
rect 10120 4410 10450 4460
rect 10900 4150 10960 4450
rect 11220 4410 11550 4460
rect 11990 4150 12050 4450
rect -6550 3300 -5420 3350
rect -4160 3300 -3870 3350
rect -2890 3300 -2480 3350
rect -1520 3300 -1110 3350
rect -120 3300 180 3350
rect 2550 3300 2850 3350
rect 3850 3300 4150 3350
rect 5250 3300 5550 3350
rect 6600 3300 6900 3350
rect 9040 3300 9370 3350
rect 10140 3300 10470 3350
rect 11190 3300 11520 3350
rect -6550 2800 -5420 2820
rect -6550 2770 -5700 2800
rect -5710 2720 -5700 2770
rect -5460 2770 -5420 2800
rect -4100 2770 -3810 2820
rect -2860 2770 -2450 2820
rect -1510 2770 -1100 2820
rect -110 2770 190 2820
rect -5460 2720 -5450 2770
rect 970 2720 980 2820
rect 1190 2720 1200 2820
rect 1750 2720 1760 2820
rect 1970 2720 1980 2820
rect 2590 2770 2890 2820
rect 3850 2770 7610 2820
rect 7940 2770 7980 2820
rect 6408 2690 7002 2696
rect 6408 2590 6420 2690
rect 6990 2590 7002 2690
rect 6408 2584 7002 2590
rect 6000 2510 7900 2520
rect 5710 2470 7900 2510
rect -810 2370 -800 2450
rect -720 2410 -710 2450
rect -720 2370 4350 2410
rect -3030 2290 4270 2320
rect -3030 1780 -2960 2290
rect 2910 2210 2920 2250
rect -1270 2180 2920 2210
rect 2990 2180 3000 2250
rect -1270 1880 -1190 2180
rect -160 2140 4160 2150
rect -170 2070 -160 2140
rect -90 2120 4160 2140
rect -90 2070 -80 2120
rect 1020 1990 1440 2060
rect -1280 1810 -1270 1880
rect -1190 1810 -1180 1880
rect 1110 1790 1120 1960
rect 1190 1790 1200 1960
rect -6340 1720 -2960 1780
rect -6340 1210 -6270 1720
rect -5490 1580 200 1660
rect -6640 1180 -6530 1210
rect -6490 1180 -6240 1210
rect -5490 1180 -5400 1580
rect -1280 1370 -1270 1440
rect -1190 1370 -1180 1440
rect -170 1370 -160 1440
rect -90 1370 -80 1440
rect -5100 1180 -1580 1210
rect -1270 1180 -1190 1370
rect -830 1270 -820 1370
rect -730 1270 -720 1370
rect -6700 690 -6670 700
rect -6460 690 -6230 700
rect -6700 670 -6230 690
rect -5100 670 -1570 700
rect -6700 -920 -6670 670
rect -4880 -410 -4850 -20
rect -4180 -410 -4150 -20
rect -5090 -440 -3650 -410
rect -3480 -440 -3450 -20
rect -6310 -480 -5720 -440
rect -6490 -920 -6480 -910
rect -6700 -950 -6480 -920
rect -6490 -970 -6480 -950
rect -6380 -970 -6370 -910
rect -6310 -950 -6280 -480
rect -6220 -670 -6210 -510
rect -6150 -670 -6140 -510
rect -6030 -670 -6020 -510
rect -5960 -670 -5950 -510
rect -5840 -670 -5830 -510
rect -5770 -670 -5760 -510
rect -6130 -910 -6120 -750
rect -6060 -910 -6050 -750
rect -5930 -910 -5920 -750
rect -5860 -910 -5850 -750
rect -5740 -910 -5730 -750
rect -5670 -910 -5660 -750
rect -5090 -950 -3650 -920
rect -6310 -990 -5810 -950
rect -820 -960 -790 1270
rect -400 1190 -390 1250
rect -240 1190 -230 1250
rect -160 1180 -90 1370
rect 120 1220 200 1580
rect 950 1560 960 1730
rect 1030 1560 1040 1730
rect 1270 1560 1280 1730
rect 1350 1560 1360 1730
rect 1390 1530 1440 1990
rect 1020 1460 1440 1530
rect 1510 1990 1930 2060
rect 4100 1990 4160 2120
rect 1510 1530 1560 1990
rect 1750 1790 1760 1960
rect 1830 1790 1840 1960
rect 4090 1930 4100 1990
rect 4160 1930 4170 1990
rect 4240 1730 4270 2290
rect 4310 1970 4350 2370
rect 5710 1980 5750 2470
rect 6050 2260 6060 2430
rect 6120 2260 6130 2430
rect 6240 2260 6250 2430
rect 6310 2260 6320 2430
rect 6440 2260 6450 2430
rect 6510 2260 6520 2430
rect 6630 2260 6640 2430
rect 6700 2260 6710 2430
rect 6820 2260 6830 2430
rect 6890 2260 6900 2430
rect 7010 2260 7020 2430
rect 7080 2260 7090 2430
rect 7200 2260 7210 2430
rect 7270 2260 7280 2430
rect 7400 2260 7410 2430
rect 7470 2260 7480 2430
rect 7590 2260 7600 2430
rect 7660 2260 7670 2430
rect 7780 2260 7790 2430
rect 7850 2260 7860 2430
rect 8190 2200 8240 2810
rect 9030 2770 9360 2820
rect 10140 2770 10470 2820
rect 11220 2770 11550 2820
rect 5960 2030 5970 2200
rect 6030 2030 6040 2200
rect 6150 2030 6160 2200
rect 6220 2030 6230 2200
rect 6340 2030 6350 2200
rect 6410 2030 6420 2200
rect 6530 2030 6540 2200
rect 6600 2030 6610 2200
rect 6720 2030 6730 2200
rect 6790 2030 6800 2200
rect 6920 2030 6930 2200
rect 6990 2030 7000 2200
rect 7110 2030 7120 2200
rect 7180 2030 7190 2200
rect 7300 2030 7310 2200
rect 7370 2030 7380 2200
rect 7490 2030 7500 2200
rect 7560 2030 7570 2200
rect 7690 2030 7700 2200
rect 7760 2030 7770 2200
rect 7880 2030 7890 2200
rect 7950 2030 7960 2200
rect 8110 2030 8120 2200
rect 8230 2030 8240 2200
rect 5710 1970 7810 1980
rect 4310 1940 7810 1970
rect 1590 1560 1600 1730
rect 1670 1560 1680 1730
rect 1910 1560 1920 1730
rect 1990 1560 2000 1730
rect 4240 1700 5670 1730
rect 2620 1590 5600 1660
rect 1510 1460 1930 1530
rect 2620 1220 2720 1590
rect 2910 1440 2920 1500
rect 2990 1440 3000 1500
rect 5570 1440 5600 1590
rect 5640 1520 5670 1700
rect 5640 1490 9090 1520
rect 120 1180 2720 1220
rect 2920 1180 2990 1440
rect 5570 1400 8280 1440
rect 4090 1310 4100 1370
rect 4160 1310 4170 1370
rect 3110 1220 3120 1250
rect 3040 1190 3120 1220
rect 3280 1190 3290 1250
rect 3040 1180 3110 1190
rect 4100 1180 4160 1310
rect 4450 1180 4770 1210
rect 4960 1180 7980 1210
rect 8210 1180 8280 1400
rect 9000 1180 9090 1490
rect 9390 1180 11890 1210
rect 4460 670 4780 700
rect 4960 670 7970 700
rect 9390 670 11890 700
rect 410 -430 440 -80
rect 570 -440 840 -410
rect 1110 -420 1140 -80
rect 1370 -440 1400 -410
rect 1390 -470 1400 -440
rect 1560 -470 1570 -410
rect 1810 -430 1840 -80
rect 1980 -440 2250 -410
rect 2510 -430 2540 -80
rect 6400 -410 6430 -40
rect 7100 -410 7130 -40
rect 6150 -440 7720 -410
rect 7800 -440 7830 -40
rect 9990 -410 10020 -80
rect 10690 -410 10720 -80
rect 11390 -410 11420 -80
rect 12090 -410 12120 -80
rect 9760 -440 12260 -410
rect -720 -770 -430 -720
rect -820 -990 -730 -960
rect -650 -980 -640 -840
rect -580 -980 -570 -840
rect -6310 -1050 -6280 -990
rect -6310 -1100 -5810 -1050
rect -6310 -1570 -6280 -1100
rect -6130 -1290 -6120 -1130
rect -6060 -1290 -6050 -1130
rect -5940 -1290 -5930 -1130
rect -5870 -1290 -5860 -1130
rect -5740 -1290 -5730 -1130
rect -5670 -1290 -5660 -1130
rect -5636 -1370 -5544 -1358
rect -6220 -1530 -6210 -1370
rect -6150 -1530 -6140 -1370
rect -6030 -1530 -6020 -1370
rect -5960 -1530 -5950 -1370
rect -5840 -1530 -5830 -1370
rect -5770 -1530 -5760 -1370
rect -5640 -1530 -5630 -1370
rect -5550 -1530 -5540 -1370
rect -820 -1460 -790 -990
rect -470 -1050 -430 -770
rect 560 -950 830 -920
rect 1290 -950 1560 -920
rect 1980 -950 2250 -920
rect 6180 -950 7750 -920
rect 9750 -950 12230 -920
rect -720 -1100 -430 -1050
rect -470 -1180 -430 -1100
rect -470 -1230 -130 -1180
rect -470 -1380 -420 -1230
rect -700 -1430 -420 -1380
rect -250 -1430 -240 -1260
rect -180 -1430 -170 -1260
rect -820 -1500 -710 -1460
rect -5636 -1542 -5544 -1530
rect -5150 -1570 -5140 -1540
rect -6310 -1600 -5140 -1570
rect -5150 -1620 -5140 -1600
rect -5050 -1570 -5040 -1540
rect -5050 -1600 -5030 -1570
rect -5050 -1620 -5040 -1600
rect -2480 -1620 -2470 -1540
rect -2370 -1590 -2360 -1540
rect -2370 -1620 -820 -1590
rect -850 -1710 -820 -1620
rect -710 -1640 -700 -1590
rect -640 -1650 -630 -1510
rect -570 -1650 -560 -1510
rect -470 -1690 -420 -1430
rect -36 -1490 46 -1478
rect -340 -1660 -330 -1490
rect -270 -1660 -260 -1490
rect -150 -1660 -140 -1490
rect -80 -1660 -70 -1490
rect -36 -1670 -30 -1490
rect 40 -1670 46 -1490
rect -36 -1682 46 -1670
rect -710 -1710 -220 -1690
rect -850 -1740 -220 -1710
<< via1 >>
rect 840 4590 1440 4750
rect 1830 4580 2310 4750
rect 1360 4400 1660 4450
rect 1360 4340 1660 4400
rect -5700 2720 -5460 2800
rect 980 2720 1190 2820
rect 1760 2720 1970 2820
rect 6420 2590 6990 2690
rect -800 2370 -720 2450
rect 2920 2180 2990 2250
rect -160 2070 -90 2140
rect -1270 1810 -1190 1880
rect 1120 1790 1190 1960
rect -1270 1370 -1190 1440
rect -160 1370 -90 1440
rect -820 1270 -730 1370
rect -6480 -970 -6380 -910
rect -6210 -670 -6150 -510
rect -6020 -670 -5960 -510
rect -5830 -670 -5770 -510
rect -6120 -910 -6060 -750
rect -5920 -910 -5860 -750
rect -5730 -910 -5670 -750
rect -390 1190 -240 1250
rect 960 1560 1030 1730
rect 1280 1560 1350 1730
rect 1760 1790 1830 1960
rect 4100 1930 4160 1990
rect 6060 2260 6120 2430
rect 6250 2260 6310 2430
rect 6450 2260 6510 2430
rect 6640 2260 6700 2430
rect 6830 2260 6890 2430
rect 7020 2260 7080 2430
rect 7210 2260 7270 2430
rect 7410 2260 7470 2430
rect 7600 2260 7660 2430
rect 7790 2260 7850 2430
rect 5970 2030 6030 2200
rect 6160 2030 6220 2200
rect 6350 2030 6410 2200
rect 6540 2030 6600 2200
rect 6730 2030 6790 2200
rect 6930 2030 6990 2200
rect 7120 2030 7180 2200
rect 7310 2030 7370 2200
rect 7500 2030 7560 2200
rect 7700 2030 7760 2200
rect 7890 2030 7950 2200
rect 8120 2030 8230 2200
rect 1600 1560 1670 1730
rect 1920 1560 1990 1730
rect 2920 1440 2990 1500
rect 4100 1310 4160 1370
rect 3120 1190 3280 1250
rect 1400 -470 1560 -410
rect -640 -980 -580 -840
rect -6120 -1290 -6060 -1130
rect -5930 -1290 -5870 -1130
rect -5730 -1290 -5670 -1130
rect -6210 -1530 -6150 -1370
rect -6020 -1530 -5960 -1370
rect -5830 -1530 -5770 -1370
rect -5630 -1530 -5550 -1370
rect -240 -1430 -180 -1260
rect -5140 -1620 -5050 -1540
rect -2470 -1620 -2370 -1540
rect -630 -1650 -570 -1510
rect -330 -1660 -270 -1490
rect -140 -1660 -80 -1490
<< metal2 >>
rect -6280 7560 -5770 7570
rect -1030 7560 -570 7580
rect -6310 7190 -6280 7560
rect -5770 7190 -1030 7560
rect -5770 7040 -5490 7190
rect -6280 7030 -5490 7040
rect -6240 5920 -5490 7030
rect -1990 6540 -1800 6550
rect -5120 6530 -1990 6540
rect -5120 6390 -5110 6530
rect -4920 6390 -1990 6530
rect -1800 6390 -1350 6540
rect -1990 6380 -1800 6390
rect -5110 6370 -4920 6380
rect -4800 6300 -4610 6310
rect -1660 6300 -1470 6310
rect -4990 6150 -4800 6300
rect -4610 6150 -1660 6300
rect -4800 6140 -4610 6150
rect -1660 6140 -1470 6150
rect -1030 5920 -570 7040
rect -6240 5550 -570 5920
rect -6240 4290 -5490 5550
rect -5110 4890 -4920 4900
rect -1990 4890 -1800 4900
rect -5120 4740 -5110 4890
rect -4920 4740 -1990 4890
rect -1800 4740 -1600 4890
rect -5110 4730 -4920 4740
rect -1990 4730 -1800 4740
rect -4800 4660 -4610 4670
rect -1660 4660 -1470 4670
rect -5000 4510 -4800 4660
rect -4610 4510 -1660 4660
rect -4800 4500 -4610 4510
rect -1660 4500 -1470 4510
rect -1030 4290 -570 5550
rect 2990 7560 3450 7580
rect 8650 7570 9100 7580
rect 8650 7560 9110 7570
rect 8470 7540 8650 7550
rect 3450 7180 8650 7540
rect 2990 5910 3450 7040
rect 8470 7040 8650 7180
rect 9110 7190 11940 7550
rect 8470 7030 9110 7040
rect 4260 6540 4450 6550
rect 4450 6530 8020 6540
rect 4450 6390 7390 6530
rect 4260 6380 4450 6390
rect 7580 6390 8020 6530
rect 7390 6370 7580 6380
rect 7700 6300 7890 6310
rect 4590 6290 4780 6300
rect 5970 6290 6190 6300
rect 4380 6140 4590 6290
rect 4780 6140 5970 6290
rect 6190 6150 7700 6290
rect 7890 6150 7900 6290
rect 6190 6140 7900 6150
rect 4590 6130 4780 6140
rect 5970 6130 6190 6140
rect 8470 5910 9100 7030
rect 9380 6540 9540 6550
rect 9370 6370 9380 6530
rect 11770 6530 11960 6540
rect 9540 6380 11770 6530
rect 9540 6370 11960 6380
rect 9380 6360 9540 6370
rect 9670 6310 9830 6320
rect 9460 6140 9670 6300
rect 12110 6300 12300 6310
rect 9830 6290 12020 6300
rect 9830 6150 10660 6290
rect 11050 6150 12020 6290
rect 9830 6140 12020 6150
rect 12110 6140 12300 6150
rect 9670 6130 9830 6140
rect 2990 5710 11920 5910
rect 2990 5550 11930 5710
rect 840 4750 1440 4760
rect 840 4580 1440 4590
rect 1830 4750 2310 4760
rect 1830 4570 2310 4580
rect 1360 4450 1660 4460
rect 1360 4330 1660 4340
rect -7240 4280 -240 4290
rect 2990 4280 3450 5550
rect 4260 4900 4450 4910
rect 4450 4890 8030 4900
rect 4450 4750 7390 4890
rect 4260 4740 4450 4750
rect 7580 4750 8030 4890
rect 7390 4730 7580 4740
rect 7700 4660 7890 4670
rect 4590 4650 4780 4660
rect 5970 4650 6190 4660
rect 4380 4500 4590 4650
rect 4780 4500 5970 4650
rect 6190 4510 7700 4650
rect 7890 4510 7900 4650
rect 6190 4500 7900 4510
rect 4590 4490 4780 4500
rect 5970 4490 6190 4500
rect 8470 4280 9100 5550
rect 9380 4900 9540 4910
rect 9370 4730 9380 4890
rect 11770 4890 11960 4900
rect 9540 4740 11770 4890
rect 9540 4730 11960 4740
rect 9380 4720 9540 4730
rect 9670 4670 9830 4680
rect 9460 4510 9670 4670
rect 9830 4660 12020 4670
rect 9830 4520 10660 4660
rect 11050 4520 12020 4660
rect 9830 4510 12020 4520
rect 12110 4660 12300 4670
rect 12110 4500 12300 4510
rect 9670 4490 9830 4500
rect -7240 4270 9100 4280
rect -7240 4080 11900 4270
rect -7240 3930 -600 4080
rect -7240 3910 -6170 3930
rect -5730 3910 -600 3930
rect -480 3910 6420 4080
rect 6990 3930 11940 4080
rect 6990 3910 8150 3930
rect 8780 3910 11940 3930
rect -600 3900 -480 3910
rect 6420 3900 6990 3910
rect -1990 3260 -1800 3270
rect 4260 3260 4450 3270
rect 9380 3260 9540 3270
rect -5110 3250 -1990 3260
rect -4920 3110 -1990 3250
rect -1800 3110 -1590 3260
rect 4450 3250 8020 3260
rect 4450 3110 7390 3250
rect -1990 3100 -1800 3110
rect 4260 3100 4450 3110
rect 7580 3110 8020 3250
rect -5110 3090 -4920 3100
rect 7390 3090 7580 3100
rect 9540 3250 12220 3260
rect 9540 3100 11770 3250
rect 11960 3100 12220 3250
rect 9540 3090 12220 3100
rect 9380 3080 9540 3090
rect 9670 3030 9830 3040
rect -4800 3020 -4610 3030
rect -1660 3020 -1470 3030
rect 7700 3020 7890 3030
rect -6870 1150 -6550 2900
rect -5700 2800 -5460 2940
rect -5700 2150 -5460 2720
rect -5000 2870 -4800 3020
rect -4610 2870 -1660 3020
rect 850 3010 1190 3020
rect 1710 3010 2050 3020
rect 4590 3010 4780 3020
rect 5970 3010 6190 3020
rect 7650 3010 7700 3020
rect -5000 2860 -4610 2870
rect -1660 2860 -1470 2870
rect -5000 2150 -4780 2860
rect -5700 1920 -4780 2150
rect -6870 1140 -6280 1150
rect -6870 980 -6600 1140
rect -6370 980 -6280 1140
rect -5700 980 -5550 1920
rect -5000 1140 -4780 1920
rect -800 2450 -720 2470
rect -1270 1880 -1190 1890
rect -1270 1440 -1190 1810
rect -800 1410 -720 2370
rect -1270 1360 -1190 1370
rect -820 1370 -720 1410
rect -820 1260 -730 1270
rect -390 1250 -240 3000
rect 1190 2860 1200 3010
rect 3130 2890 3280 3010
rect 850 2850 1190 2860
rect 1710 2850 2050 2860
rect 980 2820 1190 2850
rect -160 2140 -90 2150
rect -160 1440 -90 2070
rect 980 1960 1190 2720
rect 980 1790 1120 1960
rect 1120 1780 1190 1790
rect 1760 2820 1970 2850
rect 3100 2820 3280 2890
rect 4390 2860 4590 3010
rect 4780 2860 5970 3010
rect 6190 2870 7700 3010
rect 7890 2870 7910 3010
rect 6190 2860 7910 2870
rect 4590 2850 4780 2860
rect 5970 2850 6190 2860
rect 7650 2850 7870 2860
rect 1760 1960 1970 2720
rect 1830 1790 1970 1960
rect 1760 1780 1970 1790
rect 2920 2250 2990 2260
rect 960 1730 1030 1740
rect 1280 1730 1350 1740
rect 1600 1730 1670 1740
rect 1920 1730 1990 1740
rect 1030 1560 1280 1730
rect 1350 1560 1600 1730
rect 1670 1560 1920 1730
rect 960 1550 1990 1560
rect -160 1360 -90 1370
rect -390 1140 -240 1190
rect 1360 1140 1580 1550
rect 2920 1500 2990 2180
rect 2920 1430 2990 1440
rect 3130 1260 3280 2820
rect 6420 2690 6990 2700
rect 6420 2580 6990 2590
rect 6050 2430 7850 2440
rect 6050 2260 6060 2430
rect 6120 2260 6250 2430
rect 6310 2260 6420 2430
rect 7000 2260 7020 2430
rect 7080 2260 7210 2430
rect 7270 2260 7410 2430
rect 7470 2260 7600 2430
rect 7660 2260 7790 2430
rect 6060 2250 6120 2260
rect 6250 2250 6310 2260
rect 6420 2250 7270 2260
rect 7410 2250 7470 2260
rect 7600 2250 7660 2260
rect 7790 2250 7850 2260
rect 5970 2200 6220 2210
rect 6350 2200 6410 2210
rect 6540 2200 6600 2210
rect 6730 2200 6790 2210
rect 6930 2200 6990 2210
rect 7120 2200 7180 2210
rect 7310 2200 7370 2210
rect 7500 2200 7560 2210
rect 7700 2200 7950 2210
rect 8120 2200 8230 2210
rect 8360 2200 8550 3030
rect 9460 2860 9670 3030
rect 9830 3020 12300 3030
rect 9830 2860 10660 3020
rect 11050 2870 12110 3020
rect 11050 2860 12300 2870
rect 9470 2540 12300 2860
rect 6220 2030 6350 2200
rect 6410 2030 6540 2200
rect 6600 2030 6730 2200
rect 6790 2030 6930 2200
rect 6990 2030 7120 2200
rect 7180 2030 7310 2200
rect 7370 2030 7500 2200
rect 7560 2030 7700 2200
rect 7950 2030 8120 2200
rect 8230 2030 8550 2200
rect 6190 2020 7700 2030
rect 7900 2020 7950 2030
rect 8120 2020 8230 2030
rect 5970 2010 6190 2020
rect 7700 2010 7900 2020
rect 4100 1990 4160 2000
rect 4100 1370 4160 1930
rect 8360 1850 8550 2030
rect 4100 1300 4160 1310
rect 3120 1250 3280 1260
rect 3120 1180 3280 1190
rect 3130 1140 3280 1180
rect 5970 1140 6190 1150
rect 6810 1140 7220 1150
rect -5000 1130 -1260 1140
rect -4860 990 -3660 1130
rect -3520 990 -1260 1130
rect -5000 980 -1260 990
rect -410 980 -170 1140
rect 300 980 2640 1140
rect 3100 980 3340 1140
rect 4190 980 5970 1140
rect 6190 1130 8040 1140
rect 6190 990 6270 1130
rect 6410 990 7660 1130
rect 7880 990 8040 1130
rect 6190 980 8040 990
rect 8430 1010 8550 1850
rect 11750 1340 12300 2540
rect 9180 1150 12300 1340
rect 9180 1140 10840 1150
rect 9170 1130 10840 1140
rect 8430 980 8600 1010
rect 9170 990 9870 1130
rect 10010 990 10840 1130
rect 11230 1130 12300 1150
rect 11230 990 11870 1130
rect 12010 1050 12300 1130
rect 12010 990 12200 1050
rect 9170 980 12200 990
rect -6600 970 -6370 980
rect 5970 970 6190 980
rect 6810 970 7220 980
rect -6460 740 -6380 900
rect -5090 890 -1190 900
rect -5090 750 -4790 890
rect -4650 750 -3390 890
rect -3250 750 -1190 890
rect -5090 740 -1190 750
rect 250 740 2560 900
rect 4080 890 8040 900
rect 4080 750 6510 890
rect 6650 750 7890 890
rect 8030 750 8040 890
rect 4080 740 8040 750
rect 9090 890 12010 900
rect 9090 750 10130 890
rect 10270 750 12010 890
rect 9090 740 12010 750
rect 12160 890 12300 900
rect 12160 740 12300 750
rect -6310 100 -3010 120
rect -2780 100 -2260 120
rect -2110 100 -1560 120
rect -1410 100 5470 120
rect 5720 100 9000 120
rect -6310 90 9000 100
rect -6310 -70 12310 90
rect -6310 -240 12320 -70
rect -6180 -250 -6140 -240
rect -6600 -480 -6370 -470
rect -6620 -640 -6600 -480
rect -6370 -510 -6080 -480
rect -6020 -510 -5960 -500
rect -5830 -510 -5770 -500
rect -6370 -640 -6210 -510
rect -6600 -650 -6210 -640
rect -6480 -670 -6210 -650
rect -6150 -670 -6020 -510
rect -5960 -670 -5830 -510
rect -5770 -670 -5760 -510
rect -6480 -910 -6270 -670
rect -6210 -680 -6150 -670
rect -6020 -680 -5960 -670
rect -5830 -680 -5770 -670
rect -6120 -750 -6060 -740
rect -5920 -750 -5860 -740
rect -5730 -750 -5670 -740
rect -5620 -750 -5200 -240
rect -5000 -490 -3340 -480
rect -4860 -630 -3660 -490
rect -3520 -630 -3340 -490
rect -5000 -640 -3340 -630
rect -3050 -580 -930 -240
rect 1400 -410 1560 -400
rect -600 -540 -480 -530
rect -3050 -650 -1640 -580
rect -5040 -730 -3250 -720
rect -6170 -910 -6120 -750
rect -6060 -910 -5920 -750
rect -5860 -910 -5730 -750
rect -5670 -910 -5200 -750
rect -5090 -870 -4790 -730
rect -4650 -870 -3390 -730
rect -5090 -880 -3250 -870
rect -6380 -970 -6270 -910
rect -6120 -920 -6060 -910
rect -5920 -920 -5860 -910
rect -5730 -920 -5670 -910
rect -6480 -1130 -6270 -970
rect -6120 -1130 -6060 -1120
rect -5930 -1130 -5870 -1120
rect -5730 -1130 -5670 -1120
rect -6480 -1290 -6120 -1130
rect -6060 -1290 -5930 -1130
rect -5870 -1290 -5730 -1130
rect -5670 -1290 -5660 -1130
rect -6120 -1300 -6060 -1290
rect -5930 -1300 -5870 -1290
rect -5730 -1300 -5670 -1290
rect -5620 -1360 -5200 -910
rect -6210 -1370 -6150 -1360
rect -6020 -1370 -5960 -1360
rect -5830 -1370 -5770 -1360
rect -5630 -1370 -5200 -1360
rect -6220 -1530 -6210 -1370
rect -6150 -1530 -6020 -1370
rect -5960 -1530 -5830 -1370
rect -5770 -1530 -5630 -1370
rect -6220 -1540 -5620 -1530
rect -5660 -1860 -5620 -1540
rect -5280 -1660 -5200 -1370
rect -3050 -1020 -2060 -650
rect -1650 -670 -1640 -650
rect -600 -670 -480 -660
rect -50 -640 310 -480
rect 430 -640 2440 -470
rect -600 -830 -510 -670
rect -640 -840 -510 -830
rect -580 -930 -510 -840
rect -50 -870 130 -640
rect -640 -990 -580 -980
rect -3050 -1030 -1650 -1020
rect -3050 -1090 -2320 -1030
rect -2580 -1270 -2320 -1090
rect 200 -880 2330 -720
rect -50 -1250 130 -1230
rect -240 -1260 130 -1250
rect -180 -1430 130 -1260
rect -240 -1440 130 -1430
rect 2860 -1390 3440 -240
rect -3050 -1510 -2580 -1450
rect -330 -1490 -270 -1480
rect -140 -1490 -80 -1480
rect -5140 -1540 -5050 -1530
rect -5140 -1630 -5050 -1620
rect -4990 -1660 -2580 -1510
rect -630 -1510 -330 -1500
rect -2470 -1540 -2370 -1530
rect -2470 -1630 -2370 -1620
rect -570 -1650 -330 -1510
rect -630 -1660 -330 -1650
rect -270 -1660 -140 -1490
rect -80 -1530 200 -1490
rect -80 -1660 2860 -1530
rect -5280 -1860 -2580 -1660
rect -330 -1670 2860 -1660
rect -5620 -1870 -5280 -1860
rect 60 -1870 2860 -1670
rect 3210 -1870 3440 -1390
rect 5350 -1390 6070 -240
rect 6890 -480 7220 -470
rect 6270 -490 6890 -480
rect 6410 -630 6890 -490
rect 6270 -640 6890 -630
rect 7220 -490 7940 -480
rect 7220 -630 7660 -490
rect 7800 -630 7940 -490
rect 7220 -640 7940 -630
rect 6890 -650 7220 -640
rect 6180 -730 7850 -720
rect 6180 -870 6510 -730
rect 6650 -870 7850 -730
rect 6180 -880 7850 -870
rect 7890 -730 8030 -720
rect 7890 -880 8030 -870
rect 5350 -1840 5600 -1390
rect 2860 -1880 3210 -1870
rect 8490 -1380 9430 -240
rect 9870 -490 12220 -480
rect 10010 -630 10840 -490
rect 11230 -630 11870 -490
rect 12010 -630 12220 -490
rect 9870 -640 12220 -630
rect 9770 -730 12320 -720
rect 9770 -870 10130 -730
rect 10270 -870 12160 -730
rect 12300 -870 12320 -730
rect 9770 -880 12320 -870
rect 8490 -1530 8650 -1380
rect 6070 -1860 8650 -1530
rect 5600 -1890 6070 -1880
rect 9300 -1530 9430 -1380
rect 9300 -1550 12330 -1530
rect 9300 -1560 12350 -1550
rect 9300 -1860 11850 -1560
rect 8650 -1900 9300 -1890
rect 11850 -1900 12350 -1890
<< via2 >>
rect -6280 7040 -5770 7560
rect -1030 7040 -570 7560
rect -5110 6380 -4920 6530
rect -1990 6390 -1800 6540
rect -4800 6150 -4610 6300
rect -1660 6150 -1470 6300
rect -5110 4740 -4920 4890
rect -1990 4740 -1800 4890
rect -4800 4510 -4610 4660
rect -1660 4510 -1470 4660
rect 2990 7040 3450 7560
rect 8650 7040 9110 7560
rect 4260 6390 4450 6540
rect 7390 6380 7580 6530
rect 4590 6140 4780 6290
rect 5970 6140 6190 6290
rect 7700 6150 7890 6300
rect 9380 6370 9540 6540
rect 11770 6380 11960 6530
rect 9670 6140 9830 6310
rect 10660 6150 11050 6290
rect 12110 6150 12300 6300
rect 840 4590 1440 4750
rect 1830 4580 2310 4750
rect 1360 4340 1660 4450
rect 4260 4750 4450 4900
rect 7390 4740 7580 4890
rect 4590 4500 4780 4650
rect 5970 4500 6190 4650
rect 7700 4510 7890 4660
rect 9380 4730 9540 4900
rect 11770 4740 11960 4890
rect 9670 4500 9830 4670
rect 10660 4520 11050 4660
rect 12110 4510 12300 4660
rect -600 3910 -480 4080
rect 6420 3910 6990 4080
rect -5110 3100 -4920 3250
rect -1990 3110 -1800 3260
rect 4260 3110 4450 3260
rect 7390 3100 7580 3250
rect 9380 3090 9540 3260
rect 11770 3100 11960 3250
rect -4800 2870 -4610 3020
rect -1660 2870 -1470 3020
rect -6600 980 -6370 1140
rect 850 2860 1190 3010
rect 1710 2860 2050 3010
rect 4590 2860 4780 3010
rect 5970 2860 6190 3010
rect 7700 2870 7890 3020
rect 6420 2590 6990 2690
rect 6420 2260 6450 2430
rect 6450 2260 6510 2430
rect 6510 2260 6640 2430
rect 6640 2260 6700 2430
rect 6700 2260 6830 2430
rect 6830 2260 6890 2430
rect 6890 2260 7000 2430
rect 9670 2860 9830 3030
rect 10660 2860 11050 3020
rect 12110 2870 12300 3020
rect 5970 2030 6030 2200
rect 6030 2030 6160 2200
rect 6160 2030 6190 2200
rect 7700 2030 7760 2200
rect 7760 2030 7890 2200
rect 7890 2030 7900 2200
rect 5970 2020 6190 2030
rect 7700 2020 7900 2030
rect -5000 990 -4860 1130
rect -3660 990 -3520 1130
rect 5970 980 6190 1140
rect 6270 990 6410 1130
rect 7660 990 7880 1130
rect 9870 990 10010 1130
rect 10840 990 11230 1150
rect 11870 990 12010 1130
rect -4790 750 -4650 890
rect -3390 750 -3250 890
rect 6510 750 6650 890
rect 7890 750 8030 890
rect 10130 750 10270 890
rect 12160 750 12300 890
rect -6600 -640 -6370 -480
rect -5000 -630 -4860 -490
rect -3660 -630 -3520 -490
rect -4790 -870 -4650 -730
rect -3390 -870 -3250 -730
rect -5620 -1530 -5550 -1370
rect -5550 -1530 -5280 -1370
rect -5620 -1860 -5280 -1530
rect -2060 -1020 -1650 -650
rect -600 -660 -480 -540
rect -3050 -1450 -2580 -1090
rect -50 -1230 130 -870
rect -5140 -1620 -5050 -1540
rect -2470 -1620 -2370 -1540
rect 2860 -1870 3210 -1390
rect 6270 -630 6410 -490
rect 6890 -640 7220 -480
rect 7660 -630 7800 -490
rect 6510 -870 6650 -730
rect 7890 -870 8030 -730
rect 5600 -1880 6070 -1390
rect 9870 -630 10010 -490
rect 10840 -630 11230 -490
rect 11870 -630 12010 -490
rect 10130 -870 10270 -730
rect 12160 -870 12300 -730
rect 8650 -1890 9300 -1380
rect 11850 -1890 12350 -1560
<< metal3 >>
rect -6290 7560 -5760 7565
rect -6290 7040 -6280 7560
rect -5770 7040 -5760 7560
rect -6290 7035 -5760 7040
rect -1040 7560 -560 7565
rect -1040 7040 -1030 7560
rect -570 7040 -560 7560
rect -1040 7035 -560 7040
rect 2980 7560 3460 7565
rect 2980 7040 2990 7560
rect 3450 7040 3460 7560
rect 2980 7035 3460 7040
rect 8640 7560 9120 7565
rect 8640 7040 8650 7560
rect 9110 7040 9120 7560
rect 8640 7035 9120 7040
rect -2000 6540 -1790 6545
rect -5110 6535 -4920 6540
rect -5120 6530 -4910 6535
rect -5120 6380 -5110 6530
rect -4920 6380 -4910 6530
rect -5120 6375 -4910 6380
rect -2000 6390 -1990 6540
rect -1800 6390 -1790 6540
rect -2000 6385 -1790 6390
rect 4250 6540 4460 6545
rect 4250 6390 4260 6540
rect 4450 6390 4460 6540
rect 7390 6535 7580 6550
rect 9370 6540 9550 6545
rect 4250 6385 4460 6390
rect 7380 6530 7590 6535
rect -5110 4895 -4920 6375
rect -4800 6305 -4610 6310
rect -4810 6300 -4600 6305
rect -4810 6150 -4800 6300
rect -4610 6150 -4600 6300
rect -4810 6145 -4600 6150
rect -5120 4890 -4910 4895
rect -5120 4740 -5110 4890
rect -4920 4740 -4910 4890
rect -5120 4735 -4910 4740
rect -5110 3255 -4920 4735
rect -4800 4665 -4610 6145
rect -2000 4895 -1810 6385
rect -1670 6300 -1460 6305
rect -1670 6150 -1660 6300
rect -1470 6150 -1460 6300
rect -1670 6145 -1460 6150
rect -2000 4890 -1790 4895
rect -2000 4740 -1990 4890
rect -1800 4740 -1790 4890
rect -2000 4735 -1790 4740
rect -4810 4660 -4600 4665
rect -4810 4510 -4800 4660
rect -4610 4510 -4600 4660
rect -4810 4505 -4600 4510
rect -5120 3250 -4910 3255
rect -5120 3100 -5110 3250
rect -4920 3100 -4910 3250
rect -5120 3095 -4910 3100
rect -4800 3025 -4610 4505
rect -2000 3265 -1810 4735
rect -1660 4665 -1470 6145
rect 1800 5160 1810 5470
rect 2310 5160 2320 5470
rect 960 4755 970 4970
rect 830 4750 970 4755
rect -1670 4660 -1460 4665
rect -1670 4510 -1660 4660
rect -1470 4510 -1460 4660
rect 830 4590 840 4750
rect 830 4585 970 4590
rect -1670 4505 -1460 4510
rect 850 4540 970 4585
rect 1470 4540 1480 4970
rect 1820 4755 2290 5160
rect 4260 4905 4450 6385
rect 7380 6380 7390 6530
rect 7580 6380 7590 6530
rect 7380 6375 7590 6380
rect 4580 6290 4790 6295
rect 4580 6140 4590 6290
rect 4780 6140 4790 6290
rect 4580 6135 4790 6140
rect 5960 6290 6200 6295
rect 5960 6140 5970 6290
rect 6190 6140 6200 6290
rect 5960 6135 6200 6140
rect 4250 4900 4460 4905
rect 1820 4750 2320 4755
rect 1820 4580 1830 4750
rect 2310 4580 2320 4750
rect 4250 4750 4260 4900
rect 4450 4750 4460 4900
rect 4250 4745 4460 4750
rect 1820 4575 2320 4580
rect 1820 4570 2290 4575
rect -2000 3260 -1790 3265
rect -2000 3110 -1990 3260
rect -1800 3110 -1790 3260
rect -2000 3105 -1790 3110
rect -1660 3025 -1470 4505
rect -610 4080 -470 4085
rect -610 3910 -600 4080
rect -480 3910 -470 4080
rect -610 3905 -470 3910
rect -4810 3020 -4600 3025
rect -4810 2870 -4800 3020
rect -4610 2870 -4600 3020
rect -4810 2865 -4600 2870
rect -1670 3020 -1460 3025
rect -1670 2870 -1660 3020
rect -1470 2870 -1460 3020
rect -1670 2865 -1460 2870
rect -6610 1140 -6360 1145
rect -6610 980 -6600 1140
rect -6370 980 -6360 1140
rect -5000 1135 -4860 1140
rect -3660 1135 -3520 1140
rect -5010 1130 -4850 1135
rect -5010 990 -5000 1130
rect -4860 990 -4850 1130
rect -5010 985 -4850 990
rect -3670 1130 -3510 1135
rect -3670 990 -3660 1130
rect -3520 990 -3510 1130
rect -3670 985 -3510 990
rect -6610 -480 -6360 980
rect -6610 -640 -6600 -480
rect -6370 -640 -6360 -480
rect -5000 -485 -4860 985
rect -4790 895 -4650 900
rect -4800 890 -4640 895
rect -4800 750 -4790 890
rect -4650 750 -4640 890
rect -4800 745 -4640 750
rect -5010 -490 -4850 -485
rect -5010 -630 -5000 -490
rect -4860 -630 -4850 -490
rect -5010 -635 -4850 -630
rect -5000 -640 -4860 -635
rect -6610 -645 -6360 -640
rect -4790 -725 -4650 745
rect -3660 -485 -3520 985
rect -3390 895 -3250 900
rect -3400 890 -3240 895
rect -3400 750 -3390 890
rect -3250 750 -3240 890
rect -3400 745 -3240 750
rect -3670 -490 -3510 -485
rect -3670 -630 -3660 -490
rect -3520 -630 -3510 -490
rect -3670 -635 -3510 -630
rect -3660 -640 -3520 -635
rect -3390 -725 -3250 745
rect -600 -535 -480 3905
rect 850 3240 1200 4540
rect 1350 4450 1670 4455
rect 1350 4340 1360 4450
rect 1660 4340 1670 4450
rect 1350 4335 1670 4340
rect 4260 3265 4450 4745
rect 4590 4655 4780 6135
rect 5970 4655 6190 6135
rect 7390 4895 7580 6375
rect 9370 6370 9380 6540
rect 9540 6370 9550 6540
rect 11760 6530 11970 6535
rect 11760 6380 11770 6530
rect 11960 6380 11970 6530
rect 11760 6375 11970 6380
rect 9370 6365 9550 6370
rect 7700 6305 7890 6310
rect 7690 6300 7900 6305
rect 7690 6150 7700 6300
rect 7890 6150 7900 6300
rect 7690 6145 7900 6150
rect 7380 4890 7590 4895
rect 7380 4740 7390 4890
rect 7580 4740 7590 4890
rect 7380 4735 7590 4740
rect 4580 4650 4790 4655
rect 4580 4500 4590 4650
rect 4780 4500 4790 4650
rect 4580 4495 4790 4500
rect 5960 4650 6200 4655
rect 5960 4500 5970 4650
rect 6190 4500 6200 4650
rect 5960 4495 6200 4500
rect 4250 3260 4460 3265
rect 840 3010 1200 3240
rect 840 2860 850 3010
rect 1190 2860 1200 3010
rect 1620 3240 1850 3260
rect 1620 3030 2060 3240
rect 4250 3110 4260 3260
rect 4450 3110 4460 3260
rect 4250 3105 4460 3110
rect 1620 2860 1710 3030
rect 840 2855 1200 2860
rect 1700 2850 1710 2860
rect 2060 2850 2070 3030
rect 4590 3015 4780 4495
rect 5970 3015 6190 4495
rect 6410 4080 7000 4085
rect 6410 3910 6420 4080
rect 6990 3910 7000 4080
rect 6410 3905 7000 3910
rect 4580 3010 4790 3015
rect 4580 2860 4590 3010
rect 4780 2860 4790 3010
rect 4580 2855 4790 2860
rect 5960 3010 6200 3015
rect 5960 2860 5970 3010
rect 6190 2860 6200 3010
rect 5960 2855 6200 2860
rect 5970 2205 6190 2855
rect 6420 2695 6990 3905
rect 7390 3255 7580 4735
rect 7700 4665 7890 6145
rect 9380 4905 9540 6365
rect 9660 6310 9840 6315
rect 9660 6140 9670 6310
rect 9830 6140 9840 6310
rect 10650 6290 11060 6295
rect 10650 6150 10660 6290
rect 11050 6150 11060 6290
rect 10650 6145 11060 6150
rect 9660 6135 9840 6140
rect 9370 4900 9550 4905
rect 9370 4730 9380 4900
rect 9540 4730 9550 4900
rect 9370 4725 9550 4730
rect 7690 4660 7900 4665
rect 7690 4510 7700 4660
rect 7890 4510 7900 4660
rect 7690 4505 7900 4510
rect 7380 3250 7590 3255
rect 7380 3100 7390 3250
rect 7580 3100 7590 3250
rect 7380 3095 7590 3100
rect 7700 3040 7890 4505
rect 9380 3265 9540 4725
rect 9670 4675 9830 6135
rect 9660 4670 9840 4675
rect 9660 4500 9670 4670
rect 9830 4500 9840 4670
rect 10660 4665 11050 6145
rect 11770 4895 11960 6375
rect 12100 6300 12310 6305
rect 12100 6150 12110 6300
rect 12300 6150 12310 6300
rect 12100 6145 12310 6150
rect 11760 4890 11970 4895
rect 11760 4740 11770 4890
rect 11960 4740 11970 4890
rect 11760 4735 11970 4740
rect 10650 4660 11060 4665
rect 10650 4520 10660 4660
rect 11050 4520 11060 4660
rect 10650 4515 11060 4520
rect 9660 4495 9840 4500
rect 9370 3260 9550 3265
rect 9370 3090 9380 3260
rect 9540 3090 9550 3260
rect 9370 3085 9550 3090
rect 7700 3025 7900 3040
rect 9670 3035 9830 4495
rect 7690 3020 7900 3025
rect 7690 2870 7700 3020
rect 7890 2870 7900 3020
rect 7690 2865 7900 2870
rect 6410 2690 7000 2695
rect 6410 2590 6420 2690
rect 6990 2590 7000 2690
rect 6410 2585 7000 2590
rect 6420 2440 6990 2585
rect 6420 2435 7000 2440
rect 6410 2430 7010 2435
rect 6410 2260 6420 2430
rect 7000 2260 7010 2430
rect 6410 2255 7010 2260
rect 6740 2250 7000 2255
rect 7700 2205 7900 2865
rect 9660 3030 9840 3035
rect 9660 2860 9670 3030
rect 9830 2860 9840 3030
rect 10660 3025 11050 4515
rect 11770 3255 11960 4735
rect 12110 4665 12300 6145
rect 12100 4660 12310 4665
rect 12100 4510 12110 4660
rect 12300 4510 12310 4660
rect 12100 4505 12310 4510
rect 11760 3250 11970 3255
rect 11760 3100 11770 3250
rect 11960 3100 11970 3250
rect 11760 3095 11970 3100
rect 11770 3090 11960 3095
rect 12110 3025 12300 4505
rect 9660 2855 9840 2860
rect 10650 3020 11060 3025
rect 10650 2860 10660 3020
rect 11050 2860 11060 3020
rect 12100 3020 12310 3025
rect 12100 2870 12110 3020
rect 12300 2870 12310 3020
rect 12100 2865 12310 2870
rect 12110 2860 12300 2865
rect 10650 2855 11060 2860
rect 5960 2200 6200 2205
rect 5960 2020 5970 2200
rect 6190 2020 6200 2200
rect 5960 2015 6200 2020
rect 7690 2200 7910 2205
rect 7690 2020 7700 2200
rect 7900 2020 7910 2200
rect 7690 2015 7910 2020
rect 5970 1145 6190 2015
rect 5960 1140 6200 1145
rect 7710 1140 7890 2015
rect 10830 1150 11240 1155
rect 5960 980 5970 1140
rect 6190 1130 6430 1140
rect 7660 1135 7890 1140
rect 9870 1135 10010 1140
rect 6190 990 6270 1130
rect 6410 990 6430 1130
rect 6190 980 6430 990
rect 7650 1130 7890 1135
rect 7650 990 7660 1130
rect 7880 990 7890 1130
rect 7650 985 7890 990
rect 9860 1130 10020 1135
rect 9860 990 9870 1130
rect 10010 990 10020 1130
rect 9860 985 10020 990
rect 10830 990 10840 1150
rect 11230 990 11240 1150
rect 11870 1135 12010 1140
rect 10830 985 11240 990
rect 11860 1130 12020 1135
rect 11860 990 11870 1130
rect 12010 990 12020 1130
rect 11860 985 12020 990
rect 7660 980 7890 985
rect 5960 975 6200 980
rect 6270 -485 6410 980
rect 6510 895 6650 900
rect 6500 890 6660 895
rect 6500 750 6510 890
rect 6650 750 6660 890
rect 6500 745 6660 750
rect 6260 -490 6420 -485
rect -610 -540 -470 -535
rect -2070 -650 -1640 -645
rect -4800 -730 -4640 -725
rect -4800 -870 -4790 -730
rect -4650 -870 -4640 -730
rect -4800 -875 -4640 -870
rect -3400 -730 -3240 -725
rect -3400 -870 -3390 -730
rect -3250 -870 -3240 -730
rect -3400 -875 -3240 -870
rect -4790 -880 -4650 -875
rect -3390 -880 -3250 -875
rect -2070 -1020 -2060 -650
rect -1650 -1020 -1640 -650
rect -610 -660 -600 -540
rect -480 -660 -470 -540
rect 6260 -630 6270 -490
rect 6410 -630 6420 -490
rect 6260 -635 6420 -630
rect 6270 -640 6410 -635
rect -610 -665 -470 -660
rect 6510 -725 6650 745
rect 6890 -475 7220 960
rect 6880 -480 7230 -475
rect 6880 -640 6890 -480
rect 7220 -640 7230 -480
rect 7660 -485 7800 980
rect 7890 895 8030 900
rect 7880 890 8040 895
rect 7880 750 7890 890
rect 8030 750 8040 890
rect 7880 745 8040 750
rect 7650 -490 7810 -485
rect 7650 -630 7660 -490
rect 7800 -630 7810 -490
rect 7650 -635 7810 -630
rect 7660 -640 7800 -635
rect 6880 -645 7230 -640
rect 7890 -725 8030 745
rect 9870 -485 10010 985
rect 10130 895 10270 900
rect 10120 890 10280 895
rect 10120 750 10130 890
rect 10270 750 10280 890
rect 10120 745 10280 750
rect 9860 -490 10020 -485
rect 9860 -630 9870 -490
rect 10010 -630 10020 -490
rect 9860 -635 10020 -630
rect 9870 -640 10010 -635
rect 10130 -725 10270 745
rect 10840 -485 11230 985
rect 11870 -485 12010 985
rect 12160 895 12300 900
rect 12150 890 12310 895
rect 12150 750 12160 890
rect 12300 750 12310 890
rect 12150 745 12310 750
rect 10830 -490 11240 -485
rect 10830 -630 10840 -490
rect 11230 -630 11240 -490
rect 10830 -635 11240 -630
rect 11860 -490 12020 -485
rect 11860 -630 11870 -490
rect 12010 -630 12020 -490
rect 11860 -635 12020 -630
rect 10840 -640 11230 -635
rect 11870 -640 12010 -635
rect 12160 -725 12300 745
rect 6500 -730 6660 -725
rect -2070 -1025 -1640 -1020
rect -60 -870 140 -865
rect -3060 -1090 -2570 -1085
rect -5630 -1370 -5270 -1365
rect -5630 -1860 -5620 -1370
rect -5280 -1860 -5270 -1370
rect -3060 -1450 -3050 -1090
rect -2580 -1450 -2570 -1090
rect -3060 -1455 -2570 -1450
rect -2060 -1370 -1650 -1025
rect -60 -1230 -50 -870
rect 130 -1230 140 -870
rect 6500 -870 6510 -730
rect 6650 -870 6660 -730
rect 6500 -875 6660 -870
rect 7880 -730 8040 -725
rect 7880 -870 7890 -730
rect 8030 -870 8040 -730
rect 7880 -875 8040 -870
rect 10120 -730 10280 -725
rect 10120 -870 10130 -730
rect 10270 -870 10280 -730
rect 10120 -875 10280 -870
rect 12150 -730 12310 -725
rect 12150 -870 12160 -730
rect 12300 -870 12310 -730
rect 12150 -875 12310 -870
rect 6510 -880 6650 -875
rect 7890 -880 8030 -875
rect 10130 -880 10270 -875
rect 12160 -880 12300 -875
rect -60 -1235 140 -1230
rect -2060 -1480 -470 -1370
rect 8640 -1380 9310 -1375
rect 2850 -1390 3220 -1385
rect -5150 -1540 -5040 -1535
rect -2480 -1540 -2360 -1535
rect -5150 -1620 -5140 -1540
rect -5050 -1620 -2470 -1540
rect -2370 -1620 -2360 -1540
rect -5150 -1625 -5040 -1620
rect -2480 -1625 -2360 -1620
rect -5630 -1865 -5270 -1860
rect -2060 -1900 -900 -1480
rect -470 -1900 -460 -1480
rect 2850 -1870 2860 -1390
rect 3210 -1870 3220 -1390
rect 2850 -1875 3220 -1870
rect 5590 -1390 6080 -1385
rect 5590 -1880 5600 -1390
rect 6070 -1880 6080 -1390
rect 5590 -1885 6080 -1880
rect 8640 -1890 8650 -1380
rect 9300 -1890 9310 -1380
rect 8640 -1895 9310 -1890
rect 11840 -1560 12360 -1555
rect 11840 -1890 11850 -1560
rect 12350 -1890 12360 -1560
rect 11840 -1895 12360 -1890
<< via3 >>
rect -6280 7040 -5770 7560
rect -1030 7040 -570 7560
rect 2990 7040 3450 7560
rect 8650 7040 9110 7560
rect 1810 5160 2310 5470
rect 970 4750 1470 4970
rect 970 4590 1440 4750
rect 1440 4590 1470 4750
rect 970 4540 1470 4590
rect 1360 4340 1660 4450
rect 1710 3010 2060 3030
rect 1710 2860 2050 3010
rect 2050 2860 2060 3010
rect 1710 2850 2060 2860
rect -50 -1230 130 -870
rect -900 -1900 -470 -1480
rect 2860 -1870 3210 -1390
rect 5600 -1880 6070 -1390
rect 8650 -1890 9300 -1380
rect 11850 -1890 12350 -1560
<< metal4 >>
rect -6281 7560 -5769 7561
rect -6281 7040 -6280 7560
rect -5770 7040 -5769 7560
rect -6281 7039 -5769 7040
rect -1031 7560 -569 7561
rect -1031 7040 -1030 7560
rect -570 7040 -569 7560
rect -1031 7039 -569 7040
rect 2989 7560 3451 7561
rect 2989 7040 2990 7560
rect 3450 7040 3451 7560
rect 2989 7039 3451 7040
rect 8649 7560 9111 7561
rect 8649 7040 8650 7560
rect 9110 7040 9111 7560
rect 8649 7039 9111 7040
rect 280 5470 2360 5580
rect 280 5160 1810 5470
rect 2310 5160 2360 5470
rect 1809 5159 2311 5160
rect 969 4970 1471 4971
rect 969 4540 970 4970
rect 1470 4540 3080 4970
rect 969 4539 1471 4540
rect 1100 4450 1710 4470
rect 1100 4340 1360 4450
rect 1660 4340 1710 4450
rect 1100 4320 1710 4340
rect 1100 2470 1360 4320
rect 2060 2850 2061 3031
rect 1709 2849 2061 2850
rect -7070 -540 -6640 410
rect -51 -870 131 -869
rect -1310 -1230 -50 -870
rect 130 -1230 131 -870
rect -51 -1231 131 -1230
rect 8649 -1380 9301 -1379
rect 2859 -1390 3211 -1389
rect -901 -1480 -469 -1479
rect -901 -1900 -900 -1480
rect -470 -1900 -469 -1480
rect 2859 -1870 2860 -1390
rect 3210 -1870 3211 -1390
rect 2859 -1871 3211 -1870
rect 5599 -1390 6071 -1389
rect 5599 -1880 5600 -1390
rect 6070 -1880 6071 -1390
rect 5599 -1881 6071 -1880
rect 8649 -1890 8650 -1380
rect 9300 -1890 9301 -1380
rect 8649 -1891 9301 -1890
rect 11849 -1560 12351 -1559
rect 11849 -1890 11850 -1560
rect 12350 -1890 12351 -1560
rect 11849 -1891 12351 -1890
rect -901 -1901 -469 -1900
<< via4 >>
rect -6280 7040 -5770 7560
rect -1030 7040 -570 7560
rect 2990 7040 3450 7560
rect 8650 7040 9110 7560
rect 1700 3030 2060 3220
rect 1700 2850 1710 3030
rect 1710 2850 2060 3030
rect 1100 2020 1570 2470
rect -900 -1900 -470 -1480
rect 2860 -1870 3210 -1390
rect 5600 -1880 6070 -1390
rect 8650 -1890 9300 -1380
rect 11850 -1890 12350 -1560
<< metal5 >>
rect -6304 7570 -5746 7584
rect -3670 7570 -2990 7750
rect -1054 7570 -546 7584
rect 2966 7570 3474 7584
rect 4360 7570 5040 7750
rect 8626 7570 9134 7584
rect -6640 7560 12600 7570
rect -6640 7040 -6280 7560
rect -5770 7040 -1030 7560
rect -570 7040 2990 7560
rect 3450 7040 8650 7560
rect 9110 7040 12600 7560
rect -6304 7016 -5746 7040
rect -1054 7016 -546 7040
rect 2890 6510 3540 7040
rect 8626 7016 9134 7040
rect 9910 6550 10340 7040
rect 12040 6480 12600 7040
rect 1676 3220 2084 3244
rect -10 2850 1700 3220
rect 2060 2850 3230 3220
rect 1676 2826 2084 2850
rect 1076 2470 1594 2494
rect 1076 2020 1100 2470
rect 1570 2020 1594 2470
rect 1076 1996 1594 2020
rect -7070 -540 -6640 410
rect 1200 -1370 1540 1996
rect 9620 -1310 10050 190
rect 2836 -1370 3234 -1366
rect 5576 -1370 6094 -1366
rect 8590 -1370 10050 -1310
rect 11820 -1370 12600 170
rect -1580 -1380 12600 -1370
rect -1580 -1390 8650 -1380
rect -1580 -1480 2860 -1390
rect -1580 -1900 -900 -1480
rect -470 -1870 2860 -1480
rect 3210 -1870 5600 -1390
rect -470 -1880 5600 -1870
rect 6070 -1880 8650 -1390
rect -470 -1890 8650 -1880
rect 9300 -1560 12600 -1380
rect 9300 -1890 11850 -1560
rect 12350 -1890 12600 -1560
rect -470 -1900 12600 -1890
rect -924 -1924 -446 -1900
rect 2590 -1910 3420 -1900
rect 5576 -1904 6094 -1900
rect 8626 -1914 9324 -1900
rect 11820 -1930 12600 -1900
use currm_n  currm_n_0
timestamp 1653925904
transform 1 0 820 0 1 590
box -60 -870 658 760
use currm_n  currm_n_1
timestamp 1653925904
transform 1 0 1520 0 1 590
box -60 -870 658 760
use currm_n  currm_n_2
timestamp 1653925904
transform 1 0 2220 0 1 590
box -60 -870 658 760
use currm_n  currm_n_3
timestamp 1653925904
transform 1 0 120 0 1 590
box -60 -870 658 760
use currm_n  currm_n_4
timestamp 1653925904
transform 1 0 2920 0 1 590
box -60 -870 658 760
use currm_n  currm_n_5
timestamp 1653925904
transform 1 0 -580 0 1 590
box -60 -870 658 760
use currm_n  currm_n_6
timestamp 1653925904
transform 1 0 4010 0 1 590
box -60 -870 658 760
use currm_n  currm_n_7
timestamp 1653925904
transform 1 0 4710 0 1 590
box -60 -870 658 760
use currm_n  currm_n_8
timestamp 1653925904
transform 1 0 5410 0 1 590
box -60 -870 658 760
use currm_n  currm_n_9
timestamp 1653925904
transform 1 0 7510 0 1 590
box -60 -870 658 760
use currm_n  currm_n_10
timestamp 1653925904
transform 1 0 6810 0 1 590
box -60 -870 658 760
use currm_n  currm_n_11
timestamp 1653925904
transform 1 0 6110 0 1 590
box -60 -870 658 760
use currm_n  currm_n_12
timestamp 1653925904
transform 1 0 7510 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_13
timestamp 1653925904
transform 1 0 6810 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_14
timestamp 1653925904
transform 1 0 6110 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_15
timestamp 1653925904
transform 1 0 -5170 0 1 590
box -60 -870 658 760
use currm_n  currm_n_16
timestamp 1653925904
transform 1 0 -4470 0 1 590
box -60 -870 658 760
use currm_n  currm_n_17
timestamp 1653925904
transform 1 0 -3770 0 1 590
box -60 -870 658 760
use currm_n  currm_n_18
timestamp 1653925904
transform 1 0 -2370 0 1 590
box -60 -870 658 760
use currm_n  currm_n_19
timestamp 1653925904
transform 1 0 -3070 0 1 590
box -60 -870 658 760
use currm_n  currm_n_20
timestamp 1653925904
transform 1 0 -1670 0 1 590
box -60 -870 658 760
use currm_n  currm_n_21
timestamp 1653925904
transform 1 0 -5170 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_22
timestamp 1653925904
transform 1 0 -3770 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_23
timestamp 1653925904
transform 1 0 -4470 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_31
timestamp 1653925904
transform 1 0 -6700 0 1 590
box -60 -870 658 760
use currm_n  currm_n_32
timestamp 1653925904
transform 1 0 11800 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_33
timestamp 1653925904
transform 1 0 -5870 0 1 590
box -60 -870 658 760
use currm_n  currm_n_35
timestamp 1653925904
transform 1 0 9700 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_36
timestamp 1653925904
transform 1 0 10400 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_37
timestamp 1653925904
transform 1 0 11100 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_38
timestamp 1653925904
transform 1 0 9000 0 1 590
box -60 -870 658 760
use currm_n  currm_n_39
timestamp 1653925904
transform 1 0 11100 0 1 590
box -60 -870 658 760
use currm_n  currm_n_40
timestamp 1653925904
transform 1 0 10400 0 1 590
box -60 -870 658 760
use currm_n  currm_n_41
timestamp 1653925904
transform 1 0 9700 0 1 590
box -60 -870 658 760
use currm_n  currm_n_42
timestamp 1653925904
transform 1 0 11800 0 1 590
box -60 -870 658 760
use currm_n  currm_n_43
timestamp 1653925904
transform 1 0 8210 0 1 590
box -60 -870 658 760
use currm_n  currm_n_44
timestamp 1653925904
transform 1 0 1520 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_45
timestamp 1653925904
transform 1 0 2220 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_46
timestamp 1653925904
transform 1 0 120 0 1 -1030
box -60 -870 658 760
use currm_n  currm_n_47
timestamp 1653925904
transform 1 0 820 0 1 -1030
box -60 -870 658 760
use currm_p  currm_p_0
timestamp 1653925904
transform 1 0 170 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_1
timestamp 1653925904
transform 1 0 1510 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_2
timestamp 1653925904
transform 1 0 -1170 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_3
timestamp 1653925904
transform 1 0 -2510 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_4
timestamp 1653925904
transform 1 0 -2510 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_5
timestamp 1653925904
transform 1 0 -2510 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_6
timestamp 1653925904
transform 1 0 -3850 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_7
timestamp 1653925904
transform 1 0 -3850 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_8
timestamp 1653925904
transform 1 0 -3850 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_9
timestamp 1653925904
transform 1 0 -5190 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_10
timestamp 1653925904
transform 1 0 -5190 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_11
timestamp 1653925904
transform 1 0 -5190 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_12
timestamp 1653925904
transform 1 0 2850 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_13
timestamp 1653925904
transform 1 0 6870 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_14
timestamp 1653925904
transform 1 0 6870 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_15
timestamp 1653925904
transform 1 0 6870 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_16
timestamp 1653925904
transform 1 0 5530 0 1 3450
box -60 -810 1298 848
use currm_p  currm_p_17
timestamp 1653925904
transform 1 0 5530 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_18
timestamp 1653925904
transform 1 0 5530 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_19
timestamp 1653925904
transform 1 0 4190 0 1 6730
box -60 -810 1298 848
use currm_p  currm_p_20
timestamp 1653925904
transform 1 0 4190 0 1 5090
box -60 -810 1298 848
use currm_p  currm_p_21
timestamp 1653925904
transform 1 0 4190 0 1 3450
box -60 -810 1298 848
use currm_ps  currm_ps_0
timestamp 1653409843
transform 1 0 8200 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_1
timestamp 1653409843
transform 1 0 9290 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_2
timestamp 1653409843
transform 1 0 9290 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_3
timestamp 1653409843
transform 1 0 9290 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_4
timestamp 1653409843
transform 1 0 10380 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_5
timestamp 1653409843
transform 1 0 10380 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_6
timestamp 1653409843
transform 1 0 10380 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_7
timestamp 1653409843
transform 1 0 11470 0 1 5970
box -50 -50 1052 1608
use currm_ps  currm_ps_8
timestamp 1653409843
transform 1 0 11470 0 1 4330
box -50 -50 1052 1608
use currm_ps  currm_ps_9
timestamp 1653409843
transform 1 0 11470 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_18
timestamp 1653409843
transform 1 0 -7380 0 1 2690
box -50 -50 1052 1608
use currm_ps  currm_ps_19
timestamp 1653409843
transform 1 0 -6290 0 1 2690
box -50 -50 1052 1608
use sky130_fd_pr__cap_mim_m3_2_D7CHNQ  sky130_fd_pr__cap_mim_m3_2_D7CHNQ_0
timestamp 1654754757
transform 0 1 4241 -1 0 3443
box -1851 -1601 1873 1601
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG#4  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_2
timestamp 1653925904
transform 0 1 -2379 -1 0 3393
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_MJMGTW#0  sky130_fd_pr__cap_mim_m3_2_MJMGTW_0
timestamp 1653911185
transform 0 1 10711 -1 0 3403
box -3351 -2101 3373 2101
use sky130_fd_pr__cap_mim_m3_2_N3PKNJ  sky130_fd_pr__cap_mim_m3_2_N3PKNJ_0
timestamp 1653911185
transform 0 -1 -6819 1 0 3291
box -3351 -1101 3373 1101
use sky130_fd_pr__cap_mim_m3_2_N3PKNJ  sky130_fd_pr__cap_mim_m3_2_N3PKNJ_1
timestamp 1653911185
transform -1 0 -4547 0 -1 -1409
box -3351 -1101 3373 1101
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_0
timestamp 1653899151
transform 1 0 -669 0 1 -1560
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_9A2JGL  sky130_fd_pr__nfet_01v8_9A2JGL_1
timestamp 1653901926
transform 1 0 -5943 0 1 -1021
box -407 -719 407 719
use sky130_fd_pr__nfet_01v8_E6B2KN  sky130_fd_pr__nfet_01v8_E6B2KN_0
timestamp 1653925904
transform 1 0 1155 0 1 1760
box -325 -410 325 410
use sky130_fd_pr__nfet_01v8_E6B2KN  sky130_fd_pr__nfet_01v8_E6B2KN_1
timestamp 1653925904
transform 1 0 1795 0 1 1760
box -325 -410 325 410
use sky130_fd_pr__nfet_01v8_lvt_LH2JGW#0  sky130_fd_pr__nfet_01v8_lvt_LH2JGW_0
timestamp 1653899151
transform 1 0 -207 0 1 -1460
box -263 -410 263 410
use sky130_fd_pr__pfet_01v8_UAQRRG  sky130_fd_pr__pfet_01v8_UAQRRG_0
timestamp 1653899151
transform 1 0 -689 0 1 -911
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_VCBWSW  sky130_fd_pr__pfet_01v8_VCBWSW_0
timestamp 1653901926
transform 1 0 6957 0 1 2229
box -1127 -419 1127 419
use sky130_fd_pr__res_xhigh_po_0p69_PAXYNN  sky130_fd_pr__res_xhigh_po_0p69_PAXYNN_0
timestamp 1654754757
transform 0 -1 1635 1 0 4662
box -235 -798 235 798
<< labels >>
rlabel metal2 1440 -640 1490 -540 1 I_Bias
rlabel metal1 -490 -1740 -440 -1690 1 Disable_FB
rlabel metal2 11870 2000 12230 2390 1 Out
rlabel metal1 1310 1990 1390 2060 1 InP
rlabel metal1 1540 1990 1620 2060 1 InN
rlabel metal5 -6580 7180 -6380 7500 1 VP
rlabel metal5 3920 -1800 4130 -1540 1 VN
rlabel metal2 1010 2480 1140 2620 1 Vm16d
rlabel metal2 1800 2470 1930 2610 1 Vm14d
<< end >>
