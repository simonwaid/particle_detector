magic
tech sky130B
magscale 1 2
timestamp 1654166568
<< locali >>
rect 1440 1340 1560 2160
rect 640 750 1410 760
rect 1440 750 1550 1340
rect 640 670 2370 750
rect 1450 660 2370 670
rect 1450 430 1550 660
rect 1450 400 1560 430
rect 1460 280 1560 400
rect 1450 20 1560 280
rect 1450 -40 1550 20
rect 2270 -40 2380 -30
rect 630 -130 2380 -40
rect 630 -540 740 -130
rect 630 -700 650 -540
rect 710 -700 740 -540
rect 630 -890 740 -700
rect 2270 -540 2380 -130
rect 2270 -700 2300 -540
rect 2360 -700 2380 -540
rect 2270 -880 2380 -700
<< viali >>
rect 650 -700 710 -540
rect 2300 -700 2360 -540
<< metal1 >>
rect 750 1600 2250 2050
rect 740 870 750 1310
rect 1340 870 1350 1310
rect 1650 870 1660 1310
rect 2250 870 2260 1310
rect 644 -540 716 -528
rect 640 -700 650 -540
rect 710 -700 720 -540
rect 644 -712 716 -700
rect 800 -770 840 -220
rect 920 -270 2190 -210
rect 920 -300 960 -270
rect 900 -700 960 -300
rect 2294 -540 2366 -528
rect 2290 -700 2300 -540
rect 2360 -700 2370 -540
rect 920 -730 960 -700
rect 2294 -712 2366 -700
rect 920 -770 2190 -730
rect 940 -790 2190 -770
<< via1 >>
rect 750 870 1340 1310
rect 1660 870 2250 1310
rect 650 -700 710 -540
rect 2300 -700 2360 -540
<< metal2 >>
rect 750 1310 1340 1320
rect 1640 1310 2280 1320
rect 720 870 750 1310
rect 1340 870 1360 1310
rect 720 360 1360 870
rect 1640 870 1660 1310
rect 2250 870 2280 1310
rect 1640 360 2280 870
rect 720 180 1400 260
rect 1610 180 2290 260
rect 720 -160 2290 180
rect 860 -460 970 -300
rect 1060 -460 2180 -160
rect 650 -540 710 -530
rect 2300 -540 2360 -530
rect 710 -700 2300 -540
rect 650 -710 710 -700
rect 2300 -710 2360 -700
use currm_comp  currm_comp_0
timestamp 1654072472
transform 1 0 710 0 1 -870
box -80 -40 1670 780
use diffamp_element_nodi  diffamp_element_nodi_0
timestamp 1654072472
transform 1 0 792 0 1 -308
box 708 208 1618 1028
use diffamp_element_nodi  diffamp_element_nodi_1
timestamp 1654072472
transform 1 0 -108 0 1 -308
box 708 208 1618 1028
use sky130_fd_pr__res_xhigh_po_2p85_8K9944  sky130_fd_pr__res_xhigh_po_2p85_8K9944_0
timestamp 1654072730
transform 1 0 1951 0 1 1458
box -451 -748 451 748
use sky130_fd_pr__res_xhigh_po_2p85_8K9944  sky130_fd_pr__res_xhigh_po_2p85_8K9944_1
timestamp 1654072730
transform 1 0 1051 0 1 1458
box -451 -748 451 748
<< labels >>
rlabel via1 970 1010 1070 1180 1 Outn
rlabel metal2 860 -460 970 -300 1 bias
rlabel metal2 860 -700 970 -540 1 VN
rlabel space 650 270 700 410 1 Inp
rlabel space 2310 270 2360 410 1 Inn
rlabel via1 1800 970 2050 1180 1 OutP
rlabel metal1 1390 1690 1600 1940 1 VP
<< end >>
