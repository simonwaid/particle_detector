magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< error_p >>
rect -845 281 -787 287
rect -653 281 -595 287
rect -461 281 -403 287
rect -269 281 -211 287
rect -77 281 -19 287
rect 115 281 173 287
rect 307 281 365 287
rect 499 281 557 287
rect 691 281 749 287
rect 883 281 941 287
rect -845 247 -833 281
rect -653 247 -641 281
rect -461 247 -449 281
rect -269 247 -257 281
rect -77 247 -65 281
rect 115 247 127 281
rect 307 247 319 281
rect 499 247 511 281
rect 691 247 703 281
rect 883 247 895 281
rect -845 241 -787 247
rect -653 241 -595 247
rect -461 241 -403 247
rect -269 241 -211 247
rect -77 241 -19 247
rect 115 241 173 247
rect 307 241 365 247
rect 499 241 557 247
rect 691 241 749 247
rect 883 241 941 247
rect -941 -247 -883 -241
rect -749 -247 -691 -241
rect -557 -247 -499 -241
rect -365 -247 -307 -241
rect -173 -247 -115 -241
rect 19 -247 77 -241
rect 211 -247 269 -241
rect 403 -247 461 -241
rect 595 -247 653 -241
rect 787 -247 845 -241
rect -941 -281 -929 -247
rect -749 -281 -737 -247
rect -557 -281 -545 -247
rect -365 -281 -353 -247
rect -173 -281 -161 -247
rect 19 -281 31 -247
rect 211 -281 223 -247
rect 403 -281 415 -247
rect 595 -281 607 -247
rect 787 -281 799 -247
rect -941 -287 -883 -281
rect -749 -287 -691 -281
rect -557 -287 -499 -281
rect -365 -287 -307 -281
rect -173 -287 -115 -281
rect 19 -287 77 -281
rect 211 -287 269 -281
rect 403 -287 461 -281
rect 595 -287 653 -281
rect 787 -287 845 -281
<< nwell >>
rect -1127 -419 1127 419
<< pmos >>
rect -927 -200 -897 200
rect -831 -200 -801 200
rect -735 -200 -705 200
rect -639 -200 -609 200
rect -543 -200 -513 200
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect 513 -200 543 200
rect 609 -200 639 200
rect 705 -200 735 200
rect 801 -200 831 200
rect 897 -200 927 200
<< pdiff >>
rect -989 188 -927 200
rect -989 -188 -977 188
rect -943 -188 -927 188
rect -989 -200 -927 -188
rect -897 188 -831 200
rect -897 -188 -881 188
rect -847 -188 -831 188
rect -897 -200 -831 -188
rect -801 188 -735 200
rect -801 -188 -785 188
rect -751 -188 -735 188
rect -801 -200 -735 -188
rect -705 188 -639 200
rect -705 -188 -689 188
rect -655 -188 -639 188
rect -705 -200 -639 -188
rect -609 188 -543 200
rect -609 -188 -593 188
rect -559 -188 -543 188
rect -609 -200 -543 -188
rect -513 188 -447 200
rect -513 -188 -497 188
rect -463 -188 -447 188
rect -513 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 513 200
rect 447 -188 463 188
rect 497 -188 513 188
rect 447 -200 513 -188
rect 543 188 609 200
rect 543 -188 559 188
rect 593 -188 609 188
rect 543 -200 609 -188
rect 639 188 705 200
rect 639 -188 655 188
rect 689 -188 705 188
rect 639 -200 705 -188
rect 735 188 801 200
rect 735 -188 751 188
rect 785 -188 801 188
rect 735 -200 801 -188
rect 831 188 897 200
rect 831 -188 847 188
rect 881 -188 897 188
rect 831 -200 897 -188
rect 927 188 989 200
rect 927 -188 943 188
rect 977 -188 989 188
rect 927 -200 989 -188
<< pdiffc >>
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
<< nsubdiff >>
rect -1091 349 -995 383
rect 995 349 1091 383
rect -1091 287 -1057 349
rect 1057 287 1091 349
rect -1091 -349 -1057 -287
rect 1057 -349 1091 -287
rect -1091 -383 -995 -349
rect 995 -383 1091 -349
<< nsubdiffcont >>
rect -995 349 995 383
rect -1091 -287 -1057 287
rect 1057 -287 1091 287
rect -995 -383 995 -349
<< poly >>
rect -849 281 -783 297
rect -849 247 -833 281
rect -799 247 -783 281
rect -849 231 -783 247
rect -657 281 -591 297
rect -657 247 -641 281
rect -607 247 -591 281
rect -657 231 -591 247
rect -465 281 -399 297
rect -465 247 -449 281
rect -415 247 -399 281
rect -465 231 -399 247
rect -273 281 -207 297
rect -273 247 -257 281
rect -223 247 -207 281
rect -273 231 -207 247
rect -81 281 -15 297
rect -81 247 -65 281
rect -31 247 -15 281
rect -81 231 -15 247
rect 111 281 177 297
rect 111 247 127 281
rect 161 247 177 281
rect 111 231 177 247
rect 303 281 369 297
rect 303 247 319 281
rect 353 247 369 281
rect 303 231 369 247
rect 495 281 561 297
rect 495 247 511 281
rect 545 247 561 281
rect 495 231 561 247
rect 687 281 753 297
rect 687 247 703 281
rect 737 247 753 281
rect 687 231 753 247
rect 879 281 945 297
rect 879 247 895 281
rect 929 247 945 281
rect 879 231 945 247
rect -927 200 -897 226
rect -831 200 -801 231
rect -735 200 -705 226
rect -639 200 -609 231
rect -543 200 -513 226
rect -447 200 -417 231
rect -351 200 -321 226
rect -255 200 -225 231
rect -159 200 -129 226
rect -63 200 -33 231
rect 33 200 63 226
rect 129 200 159 231
rect 225 200 255 226
rect 321 200 351 231
rect 417 200 447 226
rect 513 200 543 231
rect 609 200 639 226
rect 705 200 735 231
rect 801 200 831 226
rect 897 200 927 231
rect -927 -231 -897 -200
rect -831 -226 -801 -200
rect -735 -231 -705 -200
rect -639 -226 -609 -200
rect -543 -231 -513 -200
rect -447 -226 -417 -200
rect -351 -231 -321 -200
rect -255 -226 -225 -200
rect -159 -231 -129 -200
rect -63 -226 -33 -200
rect 33 -231 63 -200
rect 129 -226 159 -200
rect 225 -231 255 -200
rect 321 -226 351 -200
rect 417 -231 447 -200
rect 513 -226 543 -200
rect 609 -231 639 -200
rect 705 -226 735 -200
rect 801 -231 831 -200
rect 897 -226 927 -200
rect -945 -247 -879 -231
rect -945 -281 -929 -247
rect -895 -281 -879 -247
rect -945 -297 -879 -281
rect -753 -247 -687 -231
rect -753 -281 -737 -247
rect -703 -281 -687 -247
rect -753 -297 -687 -281
rect -561 -247 -495 -231
rect -561 -281 -545 -247
rect -511 -281 -495 -247
rect -561 -297 -495 -281
rect -369 -247 -303 -231
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -369 -297 -303 -281
rect -177 -247 -111 -231
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect -177 -297 -111 -281
rect 15 -247 81 -231
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 15 -297 81 -281
rect 207 -247 273 -231
rect 207 -281 223 -247
rect 257 -281 273 -247
rect 207 -297 273 -281
rect 399 -247 465 -231
rect 399 -281 415 -247
rect 449 -281 465 -247
rect 399 -297 465 -281
rect 591 -247 657 -231
rect 591 -281 607 -247
rect 641 -281 657 -247
rect 591 -297 657 -281
rect 783 -247 849 -231
rect 783 -281 799 -247
rect 833 -281 849 -247
rect 783 -297 849 -281
<< polycont >>
rect -833 247 -799 281
rect -641 247 -607 281
rect -449 247 -415 281
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect 511 247 545 281
rect 703 247 737 281
rect 895 247 929 281
rect -929 -281 -895 -247
rect -737 -281 -703 -247
rect -545 -281 -511 -247
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
rect 415 -281 449 -247
rect 607 -281 641 -247
rect 799 -281 833 -247
<< locali >>
rect -1091 349 -995 383
rect 995 349 1091 383
rect -1091 287 -1057 349
rect 1057 287 1091 349
rect -849 247 -833 281
rect -799 247 -783 281
rect -657 247 -641 281
rect -607 247 -591 281
rect -465 247 -449 281
rect -415 247 -399 281
rect -273 247 -257 281
rect -223 247 -207 281
rect -81 247 -65 281
rect -31 247 -15 281
rect 111 247 127 281
rect 161 247 177 281
rect 303 247 319 281
rect 353 247 369 281
rect 495 247 511 281
rect 545 247 561 281
rect 687 247 703 281
rect 737 247 753 281
rect 879 247 895 281
rect 929 247 945 281
rect -977 188 -943 204
rect -977 -204 -943 -188
rect -881 188 -847 204
rect -881 -204 -847 -188
rect -785 188 -751 204
rect -785 -204 -751 -188
rect -689 188 -655 204
rect -689 -204 -655 -188
rect -593 188 -559 204
rect -593 -204 -559 -188
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect 559 188 593 204
rect 559 -204 593 -188
rect 655 188 689 204
rect 655 -204 689 -188
rect 751 188 785 204
rect 751 -204 785 -188
rect 847 188 881 204
rect 847 -204 881 -188
rect 943 188 977 204
rect 943 -204 977 -188
rect -945 -281 -929 -247
rect -895 -281 -879 -247
rect -753 -281 -737 -247
rect -703 -281 -687 -247
rect -561 -281 -545 -247
rect -511 -281 -495 -247
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 207 -281 223 -247
rect 257 -281 273 -247
rect 399 -281 415 -247
rect 449 -281 465 -247
rect 591 -281 607 -247
rect 641 -281 657 -247
rect 783 -281 799 -247
rect 833 -281 849 -247
rect -1091 -349 -1057 -287
rect 1057 -349 1091 -287
rect -1091 -383 -995 -349
rect 995 -383 1091 -349
<< viali >>
rect -833 247 -799 281
rect -641 247 -607 281
rect -449 247 -415 281
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect 511 247 545 281
rect 703 247 737 281
rect 895 247 929 281
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect -929 -281 -895 -247
rect -737 -281 -703 -247
rect -545 -281 -511 -247
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
rect 415 -281 449 -247
rect 607 -281 641 -247
rect 799 -281 833 -247
<< metal1 >>
rect -845 281 -787 287
rect -845 247 -833 281
rect -799 247 -787 281
rect -845 241 -787 247
rect -653 281 -595 287
rect -653 247 -641 281
rect -607 247 -595 281
rect -653 241 -595 247
rect -461 281 -403 287
rect -461 247 -449 281
rect -415 247 -403 281
rect -461 241 -403 247
rect -269 281 -211 287
rect -269 247 -257 281
rect -223 247 -211 281
rect -269 241 -211 247
rect -77 281 -19 287
rect -77 247 -65 281
rect -31 247 -19 281
rect -77 241 -19 247
rect 115 281 173 287
rect 115 247 127 281
rect 161 247 173 281
rect 115 241 173 247
rect 307 281 365 287
rect 307 247 319 281
rect 353 247 365 281
rect 307 241 365 247
rect 499 281 557 287
rect 499 247 511 281
rect 545 247 557 281
rect 499 241 557 247
rect 691 281 749 287
rect 691 247 703 281
rect 737 247 749 281
rect 691 241 749 247
rect 883 281 941 287
rect 883 247 895 281
rect 929 247 941 281
rect 883 241 941 247
rect -983 188 -937 200
rect -983 -188 -977 188
rect -943 -188 -937 188
rect -983 -200 -937 -188
rect -887 188 -841 200
rect -887 -188 -881 188
rect -847 -188 -841 188
rect -887 -200 -841 -188
rect -791 188 -745 200
rect -791 -188 -785 188
rect -751 -188 -745 188
rect -791 -200 -745 -188
rect -695 188 -649 200
rect -695 -188 -689 188
rect -655 -188 -649 188
rect -695 -200 -649 -188
rect -599 188 -553 200
rect -599 -188 -593 188
rect -559 -188 -553 188
rect -599 -200 -553 -188
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect 553 188 599 200
rect 553 -188 559 188
rect 593 -188 599 188
rect 553 -200 599 -188
rect 649 188 695 200
rect 649 -188 655 188
rect 689 -188 695 188
rect 649 -200 695 -188
rect 745 188 791 200
rect 745 -188 751 188
rect 785 -188 791 188
rect 745 -200 791 -188
rect 841 188 887 200
rect 841 -188 847 188
rect 881 -188 887 188
rect 841 -200 887 -188
rect 937 188 983 200
rect 937 -188 943 188
rect 977 -188 983 188
rect 937 -200 983 -188
rect -941 -247 -883 -241
rect -941 -281 -929 -247
rect -895 -281 -883 -247
rect -941 -287 -883 -281
rect -749 -247 -691 -241
rect -749 -281 -737 -247
rect -703 -281 -691 -247
rect -749 -287 -691 -281
rect -557 -247 -499 -241
rect -557 -281 -545 -247
rect -511 -281 -499 -247
rect -557 -287 -499 -281
rect -365 -247 -307 -241
rect -365 -281 -353 -247
rect -319 -281 -307 -247
rect -365 -287 -307 -281
rect -173 -247 -115 -241
rect -173 -281 -161 -247
rect -127 -281 -115 -247
rect -173 -287 -115 -281
rect 19 -247 77 -241
rect 19 -281 31 -247
rect 65 -281 77 -247
rect 19 -287 77 -281
rect 211 -247 269 -241
rect 211 -281 223 -247
rect 257 -281 269 -247
rect 211 -287 269 -281
rect 403 -247 461 -241
rect 403 -281 415 -247
rect 449 -281 461 -247
rect 403 -287 461 -281
rect 595 -247 653 -241
rect 595 -281 607 -247
rect 641 -281 653 -247
rect 595 -287 653 -281
rect 787 -247 845 -241
rect 787 -281 799 -247
rect 833 -281 845 -247
rect 787 -287 845 -281
<< properties >>
string FIXED_BBOX -1074 -366 1074 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
