* SPICE3 file created from esd-array.ext - technology: sky130A


* Top level circuit esd-array

.end

