magic
tech sky130B
magscale 1 2
timestamp 1653990785
<< error_p >>
rect -737 272 -679 278
rect -619 272 -561 278
rect -501 272 -443 278
rect -383 272 -325 278
rect -265 272 -207 278
rect -147 272 -89 278
rect -29 272 29 278
rect 89 272 147 278
rect 207 272 265 278
rect 325 272 383 278
rect 443 272 501 278
rect 561 272 619 278
rect 679 272 737 278
rect -737 238 -725 272
rect -619 238 -607 272
rect -501 238 -489 272
rect -383 238 -371 272
rect -265 238 -253 272
rect -147 238 -135 272
rect -29 238 -17 272
rect 89 238 101 272
rect 207 238 219 272
rect 325 238 337 272
rect 443 238 455 272
rect 561 238 573 272
rect 679 238 691 272
rect -737 232 -679 238
rect -619 232 -561 238
rect -501 232 -443 238
rect -383 232 -325 238
rect -265 232 -207 238
rect -147 232 -89 238
rect -29 232 29 238
rect 89 232 147 238
rect 207 232 265 238
rect 325 232 383 238
rect 443 232 501 238
rect 561 232 619 238
rect 679 232 737 238
rect -737 -238 -679 -232
rect -619 -238 -561 -232
rect -501 -238 -443 -232
rect -383 -238 -325 -232
rect -265 -238 -207 -232
rect -147 -238 -89 -232
rect -29 -238 29 -232
rect 89 -238 147 -232
rect 207 -238 265 -232
rect 325 -238 383 -232
rect 443 -238 501 -232
rect 561 -238 619 -232
rect 679 -238 737 -232
rect -737 -272 -725 -238
rect -619 -272 -607 -238
rect -501 -272 -489 -238
rect -383 -272 -371 -238
rect -265 -272 -253 -238
rect -147 -272 -135 -238
rect -29 -272 -17 -238
rect 89 -272 101 -238
rect 207 -272 219 -238
rect 325 -272 337 -238
rect 443 -272 455 -238
rect 561 -272 573 -238
rect 679 -272 691 -238
rect -737 -278 -679 -272
rect -619 -278 -561 -272
rect -501 -278 -443 -272
rect -383 -278 -325 -272
rect -265 -278 -207 -272
rect -147 -278 -89 -272
rect -29 -278 29 -272
rect 89 -278 147 -272
rect 207 -278 265 -272
rect 325 -278 383 -272
rect 443 -278 501 -272
rect 561 -278 619 -272
rect 679 -278 737 -272
<< pwell >>
rect -934 -410 934 410
<< nmoslvt >>
rect -738 -200 -678 200
rect -620 -200 -560 200
rect -502 -200 -442 200
rect -384 -200 -324 200
rect -266 -200 -206 200
rect -148 -200 -88 200
rect -30 -200 30 200
rect 88 -200 148 200
rect 206 -200 266 200
rect 324 -200 384 200
rect 442 -200 502 200
rect 560 -200 620 200
rect 678 -200 738 200
<< ndiff >>
rect -796 188 -738 200
rect -796 -188 -784 188
rect -750 -188 -738 188
rect -796 -200 -738 -188
rect -678 188 -620 200
rect -678 -188 -666 188
rect -632 -188 -620 188
rect -678 -200 -620 -188
rect -560 188 -502 200
rect -560 -188 -548 188
rect -514 -188 -502 188
rect -560 -200 -502 -188
rect -442 188 -384 200
rect -442 -188 -430 188
rect -396 -188 -384 188
rect -442 -200 -384 -188
rect -324 188 -266 200
rect -324 -188 -312 188
rect -278 -188 -266 188
rect -324 -200 -266 -188
rect -206 188 -148 200
rect -206 -188 -194 188
rect -160 -188 -148 188
rect -206 -200 -148 -188
rect -88 188 -30 200
rect -88 -188 -76 188
rect -42 -188 -30 188
rect -88 -200 -30 -188
rect 30 188 88 200
rect 30 -188 42 188
rect 76 -188 88 188
rect 30 -200 88 -188
rect 148 188 206 200
rect 148 -188 160 188
rect 194 -188 206 188
rect 148 -200 206 -188
rect 266 188 324 200
rect 266 -188 278 188
rect 312 -188 324 188
rect 266 -200 324 -188
rect 384 188 442 200
rect 384 -188 396 188
rect 430 -188 442 188
rect 384 -200 442 -188
rect 502 188 560 200
rect 502 -188 514 188
rect 548 -188 560 188
rect 502 -200 560 -188
rect 620 188 678 200
rect 620 -188 632 188
rect 666 -188 678 188
rect 620 -200 678 -188
rect 738 188 796 200
rect 738 -188 750 188
rect 784 -188 796 188
rect 738 -200 796 -188
<< ndiffc >>
rect -784 -188 -750 188
rect -666 -188 -632 188
rect -548 -188 -514 188
rect -430 -188 -396 188
rect -312 -188 -278 188
rect -194 -188 -160 188
rect -76 -188 -42 188
rect 42 -188 76 188
rect 160 -188 194 188
rect 278 -188 312 188
rect 396 -188 430 188
rect 514 -188 548 188
rect 632 -188 666 188
rect 750 -188 784 188
<< psubdiff >>
rect -898 340 -802 374
rect 802 340 898 374
rect -898 278 -864 340
rect 864 278 898 340
rect -898 -340 -864 -278
rect 864 -340 898 -278
rect -898 -374 -802 -340
rect 802 -374 898 -340
<< psubdiffcont >>
rect -802 340 802 374
rect -898 -278 -864 278
rect 864 -278 898 278
rect -802 -374 802 -340
<< poly >>
rect -741 272 -675 288
rect -741 238 -725 272
rect -691 238 -675 272
rect -741 222 -675 238
rect -623 272 -557 288
rect -623 238 -607 272
rect -573 238 -557 272
rect -623 222 -557 238
rect -505 272 -439 288
rect -505 238 -489 272
rect -455 238 -439 272
rect -505 222 -439 238
rect -387 272 -321 288
rect -387 238 -371 272
rect -337 238 -321 272
rect -387 222 -321 238
rect -269 272 -203 288
rect -269 238 -253 272
rect -219 238 -203 272
rect -269 222 -203 238
rect -151 272 -85 288
rect -151 238 -135 272
rect -101 238 -85 272
rect -151 222 -85 238
rect -33 272 33 288
rect -33 238 -17 272
rect 17 238 33 272
rect -33 222 33 238
rect 85 272 151 288
rect 85 238 101 272
rect 135 238 151 272
rect 85 222 151 238
rect 203 272 269 288
rect 203 238 219 272
rect 253 238 269 272
rect 203 222 269 238
rect 321 272 387 288
rect 321 238 337 272
rect 371 238 387 272
rect 321 222 387 238
rect 439 272 505 288
rect 439 238 455 272
rect 489 238 505 272
rect 439 222 505 238
rect 557 272 623 288
rect 557 238 573 272
rect 607 238 623 272
rect 557 222 623 238
rect 675 272 741 288
rect 675 238 691 272
rect 725 238 741 272
rect 675 222 741 238
rect -738 200 -678 222
rect -620 200 -560 222
rect -502 200 -442 222
rect -384 200 -324 222
rect -266 200 -206 222
rect -148 200 -88 222
rect -30 200 30 222
rect 88 200 148 222
rect 206 200 266 222
rect 324 200 384 222
rect 442 200 502 222
rect 560 200 620 222
rect 678 200 738 222
rect -738 -222 -678 -200
rect -620 -222 -560 -200
rect -502 -222 -442 -200
rect -384 -222 -324 -200
rect -266 -222 -206 -200
rect -148 -222 -88 -200
rect -30 -222 30 -200
rect 88 -222 148 -200
rect 206 -222 266 -200
rect 324 -222 384 -200
rect 442 -222 502 -200
rect 560 -222 620 -200
rect 678 -222 738 -200
rect -741 -238 -675 -222
rect -741 -272 -725 -238
rect -691 -272 -675 -238
rect -741 -288 -675 -272
rect -623 -238 -557 -222
rect -623 -272 -607 -238
rect -573 -272 -557 -238
rect -623 -288 -557 -272
rect -505 -238 -439 -222
rect -505 -272 -489 -238
rect -455 -272 -439 -238
rect -505 -288 -439 -272
rect -387 -238 -321 -222
rect -387 -272 -371 -238
rect -337 -272 -321 -238
rect -387 -288 -321 -272
rect -269 -238 -203 -222
rect -269 -272 -253 -238
rect -219 -272 -203 -238
rect -269 -288 -203 -272
rect -151 -238 -85 -222
rect -151 -272 -135 -238
rect -101 -272 -85 -238
rect -151 -288 -85 -272
rect -33 -238 33 -222
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
rect 85 -238 151 -222
rect 85 -272 101 -238
rect 135 -272 151 -238
rect 85 -288 151 -272
rect 203 -238 269 -222
rect 203 -272 219 -238
rect 253 -272 269 -238
rect 203 -288 269 -272
rect 321 -238 387 -222
rect 321 -272 337 -238
rect 371 -272 387 -238
rect 321 -288 387 -272
rect 439 -238 505 -222
rect 439 -272 455 -238
rect 489 -272 505 -238
rect 439 -288 505 -272
rect 557 -238 623 -222
rect 557 -272 573 -238
rect 607 -272 623 -238
rect 557 -288 623 -272
rect 675 -238 741 -222
rect 675 -272 691 -238
rect 725 -272 741 -238
rect 675 -288 741 -272
<< polycont >>
rect -725 238 -691 272
rect -607 238 -573 272
rect -489 238 -455 272
rect -371 238 -337 272
rect -253 238 -219 272
rect -135 238 -101 272
rect -17 238 17 272
rect 101 238 135 272
rect 219 238 253 272
rect 337 238 371 272
rect 455 238 489 272
rect 573 238 607 272
rect 691 238 725 272
rect -725 -272 -691 -238
rect -607 -272 -573 -238
rect -489 -272 -455 -238
rect -371 -272 -337 -238
rect -253 -272 -219 -238
rect -135 -272 -101 -238
rect -17 -272 17 -238
rect 101 -272 135 -238
rect 219 -272 253 -238
rect 337 -272 371 -238
rect 455 -272 489 -238
rect 573 -272 607 -238
rect 691 -272 725 -238
<< locali >>
rect -898 340 -802 374
rect 802 340 898 374
rect -898 278 -864 340
rect 864 278 898 340
rect -741 238 -725 272
rect -691 238 -675 272
rect -623 238 -607 272
rect -573 238 -557 272
rect -505 238 -489 272
rect -455 238 -439 272
rect -387 238 -371 272
rect -337 238 -321 272
rect -269 238 -253 272
rect -219 238 -203 272
rect -151 238 -135 272
rect -101 238 -85 272
rect -33 238 -17 272
rect 17 238 33 272
rect 85 238 101 272
rect 135 238 151 272
rect 203 238 219 272
rect 253 238 269 272
rect 321 238 337 272
rect 371 238 387 272
rect 439 238 455 272
rect 489 238 505 272
rect 557 238 573 272
rect 607 238 623 272
rect 675 238 691 272
rect 725 238 741 272
rect -784 188 -750 204
rect -784 -204 -750 -188
rect -666 188 -632 204
rect -666 -204 -632 -188
rect -548 188 -514 204
rect -548 -204 -514 -188
rect -430 188 -396 204
rect -430 -204 -396 -188
rect -312 188 -278 204
rect -312 -204 -278 -188
rect -194 188 -160 204
rect -194 -204 -160 -188
rect -76 188 -42 204
rect -76 -204 -42 -188
rect 42 188 76 204
rect 42 -204 76 -188
rect 160 188 194 204
rect 160 -204 194 -188
rect 278 188 312 204
rect 278 -204 312 -188
rect 396 188 430 204
rect 396 -204 430 -188
rect 514 188 548 204
rect 514 -204 548 -188
rect 632 188 666 204
rect 632 -204 666 -188
rect 750 188 784 204
rect 750 -204 784 -188
rect -741 -272 -725 -238
rect -691 -272 -675 -238
rect -623 -272 -607 -238
rect -573 -272 -557 -238
rect -505 -272 -489 -238
rect -455 -272 -439 -238
rect -387 -272 -371 -238
rect -337 -272 -321 -238
rect -269 -272 -253 -238
rect -219 -272 -203 -238
rect -151 -272 -135 -238
rect -101 -272 -85 -238
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 85 -272 101 -238
rect 135 -272 151 -238
rect 203 -272 219 -238
rect 253 -272 269 -238
rect 321 -272 337 -238
rect 371 -272 387 -238
rect 439 -272 455 -238
rect 489 -272 505 -238
rect 557 -272 573 -238
rect 607 -272 623 -238
rect 675 -272 691 -238
rect 725 -272 741 -238
rect -898 -340 -864 -278
rect 864 -340 898 -278
rect -898 -374 -802 -340
rect 802 -374 898 -340
<< viali >>
rect -725 238 -691 272
rect -607 238 -573 272
rect -489 238 -455 272
rect -371 238 -337 272
rect -253 238 -219 272
rect -135 238 -101 272
rect -17 238 17 272
rect 101 238 135 272
rect 219 238 253 272
rect 337 238 371 272
rect 455 238 489 272
rect 573 238 607 272
rect 691 238 725 272
rect -784 -188 -750 188
rect -666 -188 -632 188
rect -548 -188 -514 188
rect -430 -188 -396 188
rect -312 -188 -278 188
rect -194 -188 -160 188
rect -76 -188 -42 188
rect 42 -188 76 188
rect 160 -188 194 188
rect 278 -188 312 188
rect 396 -188 430 188
rect 514 -188 548 188
rect 632 -188 666 188
rect 750 -188 784 188
rect -725 -272 -691 -238
rect -607 -272 -573 -238
rect -489 -272 -455 -238
rect -371 -272 -337 -238
rect -253 -272 -219 -238
rect -135 -272 -101 -238
rect -17 -272 17 -238
rect 101 -272 135 -238
rect 219 -272 253 -238
rect 337 -272 371 -238
rect 455 -272 489 -238
rect 573 -272 607 -238
rect 691 -272 725 -238
<< metal1 >>
rect -737 272 -679 278
rect -737 238 -725 272
rect -691 238 -679 272
rect -737 232 -679 238
rect -619 272 -561 278
rect -619 238 -607 272
rect -573 238 -561 272
rect -619 232 -561 238
rect -501 272 -443 278
rect -501 238 -489 272
rect -455 238 -443 272
rect -501 232 -443 238
rect -383 272 -325 278
rect -383 238 -371 272
rect -337 238 -325 272
rect -383 232 -325 238
rect -265 272 -207 278
rect -265 238 -253 272
rect -219 238 -207 272
rect -265 232 -207 238
rect -147 272 -89 278
rect -147 238 -135 272
rect -101 238 -89 272
rect -147 232 -89 238
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect 89 272 147 278
rect 89 238 101 272
rect 135 238 147 272
rect 89 232 147 238
rect 207 272 265 278
rect 207 238 219 272
rect 253 238 265 272
rect 207 232 265 238
rect 325 272 383 278
rect 325 238 337 272
rect 371 238 383 272
rect 325 232 383 238
rect 443 272 501 278
rect 443 238 455 272
rect 489 238 501 272
rect 443 232 501 238
rect 561 272 619 278
rect 561 238 573 272
rect 607 238 619 272
rect 561 232 619 238
rect 679 272 737 278
rect 679 238 691 272
rect 725 238 737 272
rect 679 232 737 238
rect -790 188 -744 200
rect -790 -188 -784 188
rect -750 -188 -744 188
rect -790 -200 -744 -188
rect -672 188 -626 200
rect -672 -188 -666 188
rect -632 -188 -626 188
rect -672 -200 -626 -188
rect -554 188 -508 200
rect -554 -188 -548 188
rect -514 -188 -508 188
rect -554 -200 -508 -188
rect -436 188 -390 200
rect -436 -188 -430 188
rect -396 -188 -390 188
rect -436 -200 -390 -188
rect -318 188 -272 200
rect -318 -188 -312 188
rect -278 -188 -272 188
rect -318 -200 -272 -188
rect -200 188 -154 200
rect -200 -188 -194 188
rect -160 -188 -154 188
rect -200 -200 -154 -188
rect -82 188 -36 200
rect -82 -188 -76 188
rect -42 -188 -36 188
rect -82 -200 -36 -188
rect 36 188 82 200
rect 36 -188 42 188
rect 76 -188 82 188
rect 36 -200 82 -188
rect 154 188 200 200
rect 154 -188 160 188
rect 194 -188 200 188
rect 154 -200 200 -188
rect 272 188 318 200
rect 272 -188 278 188
rect 312 -188 318 188
rect 272 -200 318 -188
rect 390 188 436 200
rect 390 -188 396 188
rect 430 -188 436 188
rect 390 -200 436 -188
rect 508 188 554 200
rect 508 -188 514 188
rect 548 -188 554 188
rect 508 -200 554 -188
rect 626 188 672 200
rect 626 -188 632 188
rect 666 -188 672 188
rect 626 -200 672 -188
rect 744 188 790 200
rect 744 -188 750 188
rect 784 -188 790 188
rect 744 -200 790 -188
rect -737 -238 -679 -232
rect -737 -272 -725 -238
rect -691 -272 -679 -238
rect -737 -278 -679 -272
rect -619 -238 -561 -232
rect -619 -272 -607 -238
rect -573 -272 -561 -238
rect -619 -278 -561 -272
rect -501 -238 -443 -232
rect -501 -272 -489 -238
rect -455 -272 -443 -238
rect -501 -278 -443 -272
rect -383 -238 -325 -232
rect -383 -272 -371 -238
rect -337 -272 -325 -238
rect -383 -278 -325 -272
rect -265 -238 -207 -232
rect -265 -272 -253 -238
rect -219 -272 -207 -238
rect -265 -278 -207 -272
rect -147 -238 -89 -232
rect -147 -272 -135 -238
rect -101 -272 -89 -238
rect -147 -278 -89 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 89 -238 147 -232
rect 89 -272 101 -238
rect 135 -272 147 -238
rect 89 -278 147 -272
rect 207 -238 265 -232
rect 207 -272 219 -238
rect 253 -272 265 -238
rect 207 -278 265 -272
rect 325 -238 383 -232
rect 325 -272 337 -238
rect 371 -272 383 -238
rect 325 -278 383 -272
rect 443 -238 501 -232
rect 443 -272 455 -238
rect 489 -272 501 -238
rect 443 -278 501 -272
rect 561 -238 619 -232
rect 561 -272 573 -238
rect 607 -272 619 -238
rect 561 -278 619 -272
rect 679 -238 737 -232
rect 679 -272 691 -238
rect 725 -272 737 -238
rect 679 -278 737 -272
<< properties >>
string FIXED_BBOX -881 -357 881 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.3 m 1 nf 13 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
