magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< pwell >>
rect 82 1150 2452 1216
rect 82 640 2452 706
rect 82 532 2452 598
rect 82 22 2452 88
<< poly >>
rect 82 1200 2452 1216
rect 82 1166 194 1200
rect 228 1166 386 1200
rect 420 1166 578 1200
rect 612 1166 770 1200
rect 804 1166 962 1200
rect 996 1166 1154 1200
rect 1188 1166 1346 1200
rect 1380 1166 1538 1200
rect 1572 1166 1730 1200
rect 1764 1166 1922 1200
rect 1956 1166 2114 1200
rect 2148 1166 2306 1200
rect 2340 1166 2452 1200
rect 82 1150 2452 1166
rect 82 690 2452 706
rect 82 656 98 690
rect 132 656 290 690
rect 324 656 482 690
rect 516 656 674 690
rect 708 656 866 690
rect 900 656 1058 690
rect 1092 656 1250 690
rect 1284 656 1442 690
rect 1476 656 1634 690
rect 1668 656 1826 690
rect 1860 656 2018 690
rect 2052 656 2210 690
rect 2244 656 2402 690
rect 2436 656 2452 690
rect 82 640 2452 656
rect 82 582 2452 598
rect 82 548 98 582
rect 132 548 290 582
rect 324 548 482 582
rect 516 548 674 582
rect 708 548 866 582
rect 900 548 1058 582
rect 1092 548 1250 582
rect 1284 548 1442 582
rect 1476 548 1634 582
rect 1668 548 1826 582
rect 1860 548 2018 582
rect 2052 548 2210 582
rect 2244 548 2402 582
rect 2436 548 2452 582
rect 82 532 2452 548
rect 82 72 2452 88
rect 82 38 194 72
rect 228 38 386 72
rect 420 38 578 72
rect 612 38 770 72
rect 804 38 962 72
rect 996 38 1154 72
rect 1188 38 1346 72
rect 1380 38 1538 72
rect 1572 38 1730 72
rect 1764 38 1922 72
rect 1956 38 2114 72
rect 2148 38 2306 72
rect 2340 38 2452 72
rect 82 22 2452 38
<< polycont >>
rect 194 1166 228 1200
rect 386 1166 420 1200
rect 578 1166 612 1200
rect 770 1166 804 1200
rect 962 1166 996 1200
rect 1154 1166 1188 1200
rect 1346 1166 1380 1200
rect 1538 1166 1572 1200
rect 1730 1166 1764 1200
rect 1922 1166 1956 1200
rect 2114 1166 2148 1200
rect 2306 1166 2340 1200
rect 98 656 132 690
rect 290 656 324 690
rect 482 656 516 690
rect 674 656 708 690
rect 866 656 900 690
rect 1058 656 1092 690
rect 1250 656 1284 690
rect 1442 656 1476 690
rect 1634 656 1668 690
rect 1826 656 1860 690
rect 2018 656 2052 690
rect 2210 656 2244 690
rect 2402 656 2436 690
rect 98 548 132 582
rect 290 548 324 582
rect 482 548 516 582
rect 674 548 708 582
rect 866 548 900 582
rect 1058 548 1092 582
rect 1250 548 1284 582
rect 1442 548 1476 582
rect 1634 548 1668 582
rect 1826 548 1860 582
rect 2018 548 2052 582
rect 2210 548 2244 582
rect 2402 548 2436 582
rect 194 38 228 72
rect 386 38 420 72
rect 578 38 612 72
rect 770 38 804 72
rect 962 38 996 72
rect 1154 38 1188 72
rect 1346 38 1380 72
rect 1538 38 1572 72
rect 1730 38 1764 72
rect 1922 38 1956 72
rect 2114 38 2148 72
rect 2306 38 2340 72
<< locali >>
rect 82 1166 194 1200
rect 228 1166 386 1200
rect 420 1166 578 1200
rect 612 1166 770 1200
rect 804 1166 962 1200
rect 996 1166 1154 1200
rect 1188 1166 1346 1200
rect 1380 1166 1538 1200
rect 1572 1166 1730 1200
rect 1764 1166 1922 1200
rect 1956 1166 2114 1200
rect 2148 1166 2306 1200
rect 2340 1166 2452 1200
rect 82 656 98 690
rect 132 656 290 690
rect 324 656 482 690
rect 516 656 674 690
rect 708 656 866 690
rect 900 656 1058 690
rect 1092 656 1250 690
rect 1284 656 1442 690
rect 1476 656 1634 690
rect 1668 656 1826 690
rect 1860 656 2018 690
rect 2052 656 2210 690
rect 2244 656 2402 690
rect 2436 656 2452 690
rect 82 548 98 582
rect 132 548 290 582
rect 324 548 482 582
rect 516 548 674 582
rect 708 548 866 582
rect 900 548 1058 582
rect 1092 548 1250 582
rect 1284 548 1442 582
rect 1476 548 1634 582
rect 1668 548 1826 582
rect 1860 548 2018 582
rect 2052 548 2210 582
rect 2244 548 2402 582
rect 2436 548 2452 582
rect 82 38 194 72
rect 228 38 386 72
rect 420 38 578 72
rect 612 38 770 72
rect 804 38 962 72
rect 996 38 1154 72
rect 1188 38 1346 72
rect 1380 38 1538 72
rect 1572 38 1730 72
rect 1764 38 1922 72
rect 1956 38 2114 72
rect 2148 38 2306 72
rect 2340 38 2452 72
<< viali >>
rect 194 1166 228 1200
rect 386 1166 420 1200
rect 578 1166 612 1200
rect 770 1166 804 1200
rect 962 1166 996 1200
rect 1154 1166 1188 1200
rect 1346 1166 1380 1200
rect 1538 1166 1572 1200
rect 1730 1166 1764 1200
rect 1922 1166 1956 1200
rect 2114 1166 2148 1200
rect 2306 1166 2340 1200
rect 98 656 132 690
rect 290 656 324 690
rect 482 656 516 690
rect 674 656 708 690
rect 866 656 900 690
rect 1058 656 1092 690
rect 1250 656 1284 690
rect 1442 656 1476 690
rect 1634 656 1668 690
rect 1826 656 1860 690
rect 2018 656 2052 690
rect 2210 656 2244 690
rect 2402 656 2436 690
rect 98 548 132 582
rect 290 548 324 582
rect 482 548 516 582
rect 674 548 708 582
rect 866 548 900 582
rect 1058 548 1092 582
rect 1250 548 1284 582
rect 1442 548 1476 582
rect 1634 548 1668 582
rect 1826 548 1860 582
rect 2018 548 2052 582
rect 2210 548 2244 582
rect 2402 548 2436 582
rect 194 38 228 72
rect 386 38 420 72
rect 578 38 612 72
rect 770 38 804 72
rect 962 38 996 72
rect 1154 38 1188 72
rect 1346 38 1380 72
rect 1538 38 1572 72
rect 1730 38 1764 72
rect 1922 38 1956 72
rect 2114 38 2148 72
rect 2306 38 2340 72
<< metal1 >>
rect -10 1200 2540 1270
rect -10 1166 194 1200
rect 228 1166 386 1200
rect 420 1166 578 1200
rect 612 1166 770 1200
rect 804 1166 962 1200
rect 996 1166 1154 1200
rect 1188 1166 1346 1200
rect 1380 1166 1538 1200
rect 1572 1166 1730 1200
rect 1764 1166 1922 1200
rect 1956 1166 2114 1200
rect 2148 1166 2306 1200
rect 2340 1166 2540 1200
rect -10 1160 2540 1166
rect 126 952 136 1128
rect 190 952 200 1128
rect 318 952 328 1128
rect 382 952 392 1128
rect 510 952 520 1128
rect 574 952 584 1128
rect 702 952 712 1128
rect 766 952 776 1128
rect 894 952 904 1128
rect 958 952 968 1128
rect 1086 952 1096 1128
rect 1150 952 1160 1128
rect 1278 952 1288 1128
rect 1342 952 1352 1128
rect 1470 952 1480 1128
rect 1534 952 1544 1128
rect 1662 952 1672 1128
rect 1726 952 1736 1128
rect 1854 952 1864 1128
rect 1918 952 1928 1128
rect 2046 952 2056 1128
rect 2110 952 2120 1128
rect 2238 952 2248 1128
rect 2302 952 2312 1128
rect 2430 952 2440 1128
rect 2494 952 2504 1128
rect 30 728 40 904
rect 94 728 104 904
rect 222 728 232 904
rect 286 728 296 904
rect 414 728 424 904
rect 478 728 488 904
rect 606 728 616 904
rect 670 728 680 904
rect 798 728 808 904
rect 862 728 872 904
rect 990 728 1000 904
rect 1054 728 1064 904
rect 1182 728 1192 904
rect 1246 728 1256 904
rect 1374 728 1384 904
rect 1438 728 1448 904
rect 1566 728 1576 904
rect 1630 728 1640 904
rect 1758 728 1768 904
rect 1822 728 1832 904
rect 1950 728 1960 904
rect 2014 728 2024 904
rect 2142 728 2152 904
rect 2206 728 2216 904
rect 2334 728 2344 904
rect 2398 728 2408 904
rect -10 690 2540 700
rect -10 656 98 690
rect 132 656 290 690
rect 324 656 482 690
rect 516 656 674 690
rect 708 656 866 690
rect 900 656 1058 690
rect 1092 656 1250 690
rect 1284 656 1442 690
rect 1476 656 1634 690
rect 1668 656 1826 690
rect 1860 656 2018 690
rect 2052 656 2210 690
rect 2244 656 2402 690
rect 2436 656 2540 690
rect -10 582 2540 656
rect -10 548 98 582
rect 132 548 290 582
rect 324 548 482 582
rect 516 548 674 582
rect 708 548 866 582
rect 900 548 1058 582
rect 1092 548 1250 582
rect 1284 548 1442 582
rect 1476 548 1634 582
rect 1668 548 1826 582
rect 1860 548 2018 582
rect 2052 548 2210 582
rect 2244 548 2402 582
rect 2436 548 2540 582
rect -10 540 2540 548
rect 126 334 136 510
rect 190 334 200 510
rect 318 334 328 510
rect 382 334 392 510
rect 510 334 520 510
rect 574 334 584 510
rect 702 334 712 510
rect 766 334 776 510
rect 894 334 904 510
rect 958 334 968 510
rect 1086 334 1096 510
rect 1150 334 1160 510
rect 1278 334 1288 510
rect 1342 334 1352 510
rect 1470 334 1480 510
rect 1534 334 1544 510
rect 1662 334 1672 510
rect 1726 334 1736 510
rect 1854 334 1864 510
rect 1918 334 1928 510
rect 2046 334 2056 510
rect 2110 334 2120 510
rect 2238 334 2248 510
rect 2302 334 2312 510
rect 2430 334 2440 510
rect 2494 334 2504 510
rect 30 110 40 286
rect 94 110 104 286
rect 222 110 232 286
rect 286 110 296 286
rect 414 110 424 286
rect 478 110 488 286
rect 606 110 616 286
rect 670 110 680 286
rect 798 110 808 286
rect 862 110 872 286
rect 990 110 1000 286
rect 1054 110 1064 286
rect 1182 110 1192 286
rect 1246 110 1256 286
rect 1374 110 1384 286
rect 1438 110 1448 286
rect 1566 110 1576 286
rect 1630 110 1640 286
rect 1758 110 1768 286
rect 1822 110 1832 286
rect 1950 110 1960 286
rect 2014 110 2024 286
rect 2142 110 2152 286
rect 2206 110 2216 286
rect 2334 110 2344 286
rect 2398 110 2408 286
rect -10 72 2540 80
rect -10 38 194 72
rect 228 38 386 72
rect 420 38 578 72
rect 612 38 770 72
rect 804 38 962 72
rect 996 38 1154 72
rect 1188 38 1346 72
rect 1380 38 1538 72
rect 1572 38 1730 72
rect 1764 38 1922 72
rect 1956 38 2114 72
rect 2148 38 2306 72
rect 2340 38 2540 72
rect -10 -30 2540 38
<< via1 >>
rect 136 952 190 1128
rect 328 952 382 1128
rect 520 952 574 1128
rect 712 952 766 1128
rect 904 952 958 1128
rect 1096 952 1150 1128
rect 1288 952 1342 1128
rect 1480 952 1534 1128
rect 1672 952 1726 1128
rect 1864 952 1918 1128
rect 2056 952 2110 1128
rect 2248 952 2302 1128
rect 2440 952 2494 1128
rect 40 728 94 904
rect 232 728 286 904
rect 424 728 478 904
rect 616 728 670 904
rect 808 728 862 904
rect 1000 728 1054 904
rect 1192 728 1246 904
rect 1384 728 1438 904
rect 1576 728 1630 904
rect 1768 728 1822 904
rect 1960 728 2014 904
rect 2152 728 2206 904
rect 2344 728 2398 904
rect 136 334 190 510
rect 328 334 382 510
rect 520 334 574 510
rect 712 334 766 510
rect 904 334 958 510
rect 1096 334 1150 510
rect 1288 334 1342 510
rect 1480 334 1534 510
rect 1672 334 1726 510
rect 1864 334 1918 510
rect 2056 334 2110 510
rect 2248 334 2302 510
rect 2440 334 2494 510
rect 40 110 94 286
rect 232 110 286 286
rect 424 110 478 286
rect 616 110 670 286
rect 808 110 862 286
rect 1000 110 1054 286
rect 1192 110 1246 286
rect 1384 110 1438 286
rect 1576 110 1630 286
rect 1768 110 1822 286
rect 1960 110 2014 286
rect 2152 110 2206 286
rect 2344 110 2398 286
<< metal2 >>
rect 30 1128 2500 1140
rect 30 980 136 1128
rect 190 980 328 1128
rect 136 942 190 952
rect 382 980 520 1128
rect 328 942 382 952
rect 574 980 712 1128
rect 520 942 574 952
rect 766 980 904 1128
rect 712 942 766 952
rect 958 980 1096 1128
rect 904 942 958 952
rect 1150 980 1288 1128
rect 1096 942 1150 952
rect 1342 980 1480 1128
rect 1288 942 1342 952
rect 1534 980 1672 1128
rect 1480 942 1534 952
rect 1726 980 1864 1128
rect 1672 942 1726 952
rect 1918 980 2056 1128
rect 1864 942 1918 952
rect 2110 980 2248 1128
rect 2056 942 2110 952
rect 2302 980 2440 1128
rect 2248 942 2302 952
rect 2494 980 2500 1128
rect 2440 942 2494 952
rect 40 904 94 914
rect 30 728 40 870
rect 232 904 286 914
rect 94 728 232 870
rect 424 904 478 914
rect 286 728 424 870
rect 616 904 670 914
rect 478 728 616 870
rect 808 904 862 914
rect 670 728 808 870
rect 1000 904 1054 914
rect 862 728 1000 870
rect 1192 904 1246 914
rect 1054 728 1192 870
rect 1384 904 1438 914
rect 1246 728 1384 870
rect 1576 904 1630 914
rect 1438 728 1576 870
rect 1768 904 1822 914
rect 1630 728 1768 870
rect 1960 904 2014 914
rect 1822 728 1960 870
rect 2152 904 2206 914
rect 2014 728 2152 870
rect 2344 904 2398 914
rect 2206 728 2344 870
rect 2398 728 2500 870
rect 30 510 2500 728
rect 30 350 136 510
rect 190 350 328 510
rect 136 324 190 334
rect 382 350 520 510
rect 328 324 382 334
rect 574 350 712 510
rect 520 324 574 334
rect 766 350 904 510
rect 712 324 766 334
rect 958 350 1096 510
rect 904 324 958 334
rect 1150 350 1288 510
rect 1096 324 1150 334
rect 1342 350 1480 510
rect 1288 324 1342 334
rect 1534 350 1672 510
rect 1480 324 1534 334
rect 1726 350 1864 510
rect 1672 324 1726 334
rect 1918 350 2056 510
rect 1864 324 1918 334
rect 2110 350 2248 510
rect 2056 324 2110 334
rect 2302 350 2440 510
rect 2248 324 2302 334
rect 2494 350 2500 510
rect 2440 324 2494 334
rect 40 286 94 296
rect 232 286 286 296
rect 94 110 232 260
rect 424 286 478 296
rect 286 110 424 260
rect 616 286 670 296
rect 478 110 616 260
rect 808 286 862 296
rect 670 110 808 260
rect 1000 286 1054 296
rect 862 110 1000 260
rect 1192 286 1246 296
rect 1054 110 1192 260
rect 1384 286 1438 296
rect 1246 110 1384 260
rect 1576 286 1630 296
rect 1438 110 1576 260
rect 1768 286 1822 296
rect 1630 110 1768 260
rect 1960 286 2014 296
rect 1822 110 1960 260
rect 2152 286 2206 296
rect 2014 110 2152 260
rect 2344 286 2398 296
rect 2206 110 2344 260
rect 2398 110 2510 260
rect 40 100 2510 110
use sky130_fd_pr__nfet_01v8_lvt_RE4MKQ  sky130_fd_pr__nfet_01v8_lvt_RE4MKQ_0
timestamp 1654760956
transform 1 0 1267 0 1 619
box -1367 -719 1367 719
<< end >>
