magic
tech sky130A
magscale 1 2
timestamp 1645542524
<< error_p >>
rect -1290 291 -230 318
rect 230 291 1290 318
rect -1290 -318 -230 -291
rect 230 -318 1290 -291
<< nwell >>
rect -1393 -291 -127 291
rect 127 -291 1393 291
<< pwell >>
rect -1503 291 1503 401
rect -1503 -291 -1393 291
rect -127 -291 127 291
rect 1393 -291 1503 291
rect -1503 -401 1503 -291
<< varactor >>
rect -1260 -200 -260 200
rect 260 -200 1260 200
<< psubdiff >>
rect -1467 331 -1371 365
rect 1371 331 1467 365
rect -1467 269 -1433 331
rect 1433 269 1467 331
rect -1467 -331 -1433 -269
rect 1433 -331 1467 -269
rect -1467 -365 -1371 -331
rect 1371 -365 1467 -331
<< nsubdiff >>
rect -1357 176 -1260 200
rect -1357 -176 -1345 176
rect -1311 -176 -1260 176
rect -1357 -200 -1260 -176
rect -260 176 -163 200
rect -260 -176 -209 176
rect -175 -176 -163 176
rect -260 -200 -163 -176
rect 163 176 260 200
rect 163 -176 175 176
rect 209 -176 260 176
rect 163 -200 260 -176
rect 1260 176 1357 200
rect 1260 -176 1311 176
rect 1345 -176 1357 176
rect 1260 -200 1357 -176
<< psubdiffcont >>
rect -1371 331 1371 365
rect -1467 -269 -1433 269
rect 1433 -269 1467 269
rect -1371 -365 1371 -331
<< nsubdiffcont >>
rect -1345 -176 -1311 176
rect -209 -176 -175 176
rect 175 -176 209 176
rect 1311 -176 1345 176
<< poly >>
rect -1260 272 -260 288
rect -1260 238 -1244 272
rect -276 238 -260 272
rect -1260 200 -260 238
rect 260 272 1260 288
rect 260 238 276 272
rect 1244 238 1260 272
rect 260 200 1260 238
rect -1260 -238 -260 -200
rect -1260 -272 -1244 -238
rect -276 -272 -260 -238
rect -1260 -288 -260 -272
rect 260 -238 1260 -200
rect 260 -272 276 -238
rect 1244 -272 1260 -238
rect 260 -288 1260 -272
<< polycont >>
rect -1244 238 -276 272
rect 276 238 1244 272
rect -1244 -272 -276 -238
rect 276 -272 1244 -238
<< locali >>
rect -1467 331 -1371 365
rect 1371 331 1467 365
rect -1467 269 -1433 331
rect -1260 238 -1244 272
rect -276 238 -260 272
rect 260 238 276 272
rect 1244 238 1260 272
rect 1433 269 1467 331
rect -1345 176 -1311 192
rect -1345 -192 -1311 -176
rect -209 176 -175 192
rect -209 -192 -175 -176
rect 175 176 209 192
rect 175 -192 209 -176
rect 1311 176 1345 192
rect 1311 -192 1345 -176
rect -1467 -331 -1433 -269
rect -1260 -272 -1244 -238
rect -276 -272 -260 -238
rect 260 -272 276 -238
rect 1244 -272 1260 -238
rect 1433 -331 1467 -269
rect -1467 -365 -1371 -331
rect 1371 -365 1467 -331
<< viali >>
rect -1244 238 -276 272
rect 276 238 1244 272
rect -1345 -176 -1311 176
rect -209 -176 -175 176
rect 175 -176 209 176
rect 1311 -176 1345 176
rect -1244 -272 -276 -238
rect 276 -272 1244 -238
<< metal1 >>
rect -1256 272 -264 278
rect -1256 238 -1244 272
rect -276 238 -264 272
rect -1256 232 -264 238
rect 264 272 1256 278
rect 264 238 276 272
rect 1244 238 1256 272
rect 264 232 1256 238
rect -1351 176 -1305 188
rect -1351 -176 -1345 176
rect -1311 -176 -1305 176
rect -1351 -188 -1305 -176
rect -215 176 -169 188
rect -215 -176 -209 176
rect -175 -176 -169 176
rect -215 -188 -169 -176
rect 169 176 215 188
rect 169 -176 175 176
rect 209 -176 215 176
rect 169 -188 215 -176
rect 1305 176 1351 188
rect 1305 -176 1311 176
rect 1345 -176 1351 176
rect 1305 -188 1351 -176
rect -1256 -238 -264 -232
rect -1256 -272 -1244 -238
rect -276 -272 -264 -238
rect -1256 -278 -264 -272
rect 264 -238 1256 -232
rect 264 -272 276 -238
rect 1244 -272 1256 -238
rect 264 -278 1256 -272
<< properties >>
string FIXED_BBOX -1450 -348 1450 348
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 2 l 5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
