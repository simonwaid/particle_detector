magic
tech sky130A
magscale 1 2
timestamp 1645787783
<< error_p >>
rect -617 281 -559 287
rect -421 281 -363 287
rect -225 281 -167 287
rect -29 281 29 287
rect 167 281 225 287
rect 363 281 421 287
rect 559 281 617 287
rect -617 247 -605 281
rect -421 247 -409 281
rect -225 247 -213 281
rect -29 247 -17 281
rect 167 247 179 281
rect 363 247 375 281
rect 559 247 571 281
rect -617 241 -559 247
rect -421 241 -363 247
rect -225 241 -167 247
rect -29 241 29 247
rect 167 241 225 247
rect 363 241 421 247
rect 559 241 617 247
rect -715 -247 -657 -241
rect -519 -247 -461 -241
rect -323 -247 -265 -241
rect -127 -247 -69 -241
rect 69 -247 127 -241
rect 265 -247 323 -241
rect 461 -247 519 -241
rect 657 -247 715 -241
rect -715 -281 -703 -247
rect -519 -281 -507 -247
rect -323 -281 -311 -247
rect -127 -281 -115 -247
rect 69 -281 81 -247
rect 265 -281 277 -247
rect 461 -281 473 -247
rect 657 -281 669 -247
rect -715 -287 -657 -281
rect -519 -287 -461 -281
rect -323 -287 -265 -281
rect -127 -287 -69 -281
rect 69 -287 127 -281
rect 265 -287 323 -281
rect 461 -287 519 -281
rect 657 -287 715 -281
<< nwell >>
rect -902 -419 902 419
<< pmos >>
rect -706 -200 -666 200
rect -608 -200 -568 200
rect -510 -200 -470 200
rect -412 -200 -372 200
rect -314 -200 -274 200
rect -216 -200 -176 200
rect -118 -200 -78 200
rect -20 -200 20 200
rect 78 -200 118 200
rect 176 -200 216 200
rect 274 -200 314 200
rect 372 -200 412 200
rect 470 -200 510 200
rect 568 -200 608 200
rect 666 -200 706 200
<< pdiff >>
rect -764 188 -706 200
rect -764 -188 -752 188
rect -718 -188 -706 188
rect -764 -200 -706 -188
rect -666 188 -608 200
rect -666 -188 -654 188
rect -620 -188 -608 188
rect -666 -200 -608 -188
rect -568 188 -510 200
rect -568 -188 -556 188
rect -522 -188 -510 188
rect -568 -200 -510 -188
rect -470 188 -412 200
rect -470 -188 -458 188
rect -424 -188 -412 188
rect -470 -200 -412 -188
rect -372 188 -314 200
rect -372 -188 -360 188
rect -326 -188 -314 188
rect -372 -200 -314 -188
rect -274 188 -216 200
rect -274 -188 -262 188
rect -228 -188 -216 188
rect -274 -200 -216 -188
rect -176 188 -118 200
rect -176 -188 -164 188
rect -130 -188 -118 188
rect -176 -200 -118 -188
rect -78 188 -20 200
rect -78 -188 -66 188
rect -32 -188 -20 188
rect -78 -200 -20 -188
rect 20 188 78 200
rect 20 -188 32 188
rect 66 -188 78 188
rect 20 -200 78 -188
rect 118 188 176 200
rect 118 -188 130 188
rect 164 -188 176 188
rect 118 -200 176 -188
rect 216 188 274 200
rect 216 -188 228 188
rect 262 -188 274 188
rect 216 -200 274 -188
rect 314 188 372 200
rect 314 -188 326 188
rect 360 -188 372 188
rect 314 -200 372 -188
rect 412 188 470 200
rect 412 -188 424 188
rect 458 -188 470 188
rect 412 -200 470 -188
rect 510 188 568 200
rect 510 -188 522 188
rect 556 -188 568 188
rect 510 -200 568 -188
rect 608 188 666 200
rect 608 -188 620 188
rect 654 -188 666 188
rect 608 -200 666 -188
rect 706 188 764 200
rect 706 -188 718 188
rect 752 -188 764 188
rect 706 -200 764 -188
<< pdiffc >>
rect -752 -188 -718 188
rect -654 -188 -620 188
rect -556 -188 -522 188
rect -458 -188 -424 188
rect -360 -188 -326 188
rect -262 -188 -228 188
rect -164 -188 -130 188
rect -66 -188 -32 188
rect 32 -188 66 188
rect 130 -188 164 188
rect 228 -188 262 188
rect 326 -188 360 188
rect 424 -188 458 188
rect 522 -188 556 188
rect 620 -188 654 188
rect 718 -188 752 188
<< nsubdiff >>
rect -866 349 -770 383
rect 770 349 866 383
rect -866 287 -832 349
rect 832 287 866 349
rect -866 -349 -832 -287
rect 832 -349 866 -287
rect -866 -383 -770 -349
rect 770 -383 866 -349
<< nsubdiffcont >>
rect -770 349 770 383
rect -866 -287 -832 287
rect 832 -287 866 287
rect -770 -383 770 -349
<< poly >>
rect -621 281 -555 297
rect -621 247 -605 281
rect -571 247 -555 281
rect -621 231 -555 247
rect -425 281 -359 297
rect -425 247 -409 281
rect -375 247 -359 281
rect -425 231 -359 247
rect -229 281 -163 297
rect -229 247 -213 281
rect -179 247 -163 281
rect -229 231 -163 247
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect 163 281 229 297
rect 163 247 179 281
rect 213 247 229 281
rect 163 231 229 247
rect 359 281 425 297
rect 359 247 375 281
rect 409 247 425 281
rect 359 231 425 247
rect 555 281 621 297
rect 555 247 571 281
rect 605 247 621 281
rect 555 231 621 247
rect -706 200 -666 226
rect -608 200 -568 231
rect -510 200 -470 226
rect -412 200 -372 231
rect -314 200 -274 226
rect -216 200 -176 231
rect -118 200 -78 226
rect -20 200 20 231
rect 78 200 118 226
rect 176 200 216 231
rect 274 200 314 226
rect 372 200 412 231
rect 470 200 510 226
rect 568 200 608 231
rect 666 200 706 226
rect -706 -231 -666 -200
rect -608 -226 -568 -200
rect -510 -231 -470 -200
rect -412 -226 -372 -200
rect -314 -231 -274 -200
rect -216 -226 -176 -200
rect -118 -231 -78 -200
rect -20 -226 20 -200
rect 78 -231 118 -200
rect 176 -226 216 -200
rect 274 -231 314 -200
rect 372 -226 412 -200
rect 470 -231 510 -200
rect 568 -226 608 -200
rect 666 -231 706 -200
rect -719 -247 -653 -231
rect -719 -281 -703 -247
rect -669 -281 -653 -247
rect -719 -297 -653 -281
rect -523 -247 -457 -231
rect -523 -281 -507 -247
rect -473 -281 -457 -247
rect -523 -297 -457 -281
rect -327 -247 -261 -231
rect -327 -281 -311 -247
rect -277 -281 -261 -247
rect -327 -297 -261 -281
rect -131 -247 -65 -231
rect -131 -281 -115 -247
rect -81 -281 -65 -247
rect -131 -297 -65 -281
rect 65 -247 131 -231
rect 65 -281 81 -247
rect 115 -281 131 -247
rect 65 -297 131 -281
rect 261 -247 327 -231
rect 261 -281 277 -247
rect 311 -281 327 -247
rect 261 -297 327 -281
rect 457 -247 523 -231
rect 457 -281 473 -247
rect 507 -281 523 -247
rect 457 -297 523 -281
rect 653 -247 719 -231
rect 653 -281 669 -247
rect 703 -281 719 -247
rect 653 -297 719 -281
<< polycont >>
rect -605 247 -571 281
rect -409 247 -375 281
rect -213 247 -179 281
rect -17 247 17 281
rect 179 247 213 281
rect 375 247 409 281
rect 571 247 605 281
rect -703 -281 -669 -247
rect -507 -281 -473 -247
rect -311 -281 -277 -247
rect -115 -281 -81 -247
rect 81 -281 115 -247
rect 277 -281 311 -247
rect 473 -281 507 -247
rect 669 -281 703 -247
<< locali >>
rect -866 349 -770 383
rect 770 349 866 383
rect -866 287 -832 349
rect 832 287 866 349
rect -621 247 -605 281
rect -571 247 -555 281
rect -425 247 -409 281
rect -375 247 -359 281
rect -229 247 -213 281
rect -179 247 -163 281
rect -33 247 -17 281
rect 17 247 33 281
rect 163 247 179 281
rect 213 247 229 281
rect 359 247 375 281
rect 409 247 425 281
rect 555 247 571 281
rect 605 247 621 281
rect -752 188 -718 204
rect -752 -204 -718 -188
rect -654 188 -620 204
rect -654 -204 -620 -188
rect -556 188 -522 204
rect -556 -204 -522 -188
rect -458 188 -424 204
rect -458 -204 -424 -188
rect -360 188 -326 204
rect -360 -204 -326 -188
rect -262 188 -228 204
rect -262 -204 -228 -188
rect -164 188 -130 204
rect -164 -204 -130 -188
rect -66 188 -32 204
rect -66 -204 -32 -188
rect 32 188 66 204
rect 32 -204 66 -188
rect 130 188 164 204
rect 130 -204 164 -188
rect 228 188 262 204
rect 228 -204 262 -188
rect 326 188 360 204
rect 326 -204 360 -188
rect 424 188 458 204
rect 424 -204 458 -188
rect 522 188 556 204
rect 522 -204 556 -188
rect 620 188 654 204
rect 620 -204 654 -188
rect 718 188 752 204
rect 718 -204 752 -188
rect -719 -281 -703 -247
rect -669 -281 -653 -247
rect -523 -281 -507 -247
rect -473 -281 -457 -247
rect -327 -281 -311 -247
rect -277 -281 -261 -247
rect -131 -281 -115 -247
rect -81 -281 -65 -247
rect 65 -281 81 -247
rect 115 -281 131 -247
rect 261 -281 277 -247
rect 311 -281 327 -247
rect 457 -281 473 -247
rect 507 -281 523 -247
rect 653 -281 669 -247
rect 703 -281 719 -247
rect -866 -349 -832 -287
rect 832 -349 866 -287
rect -866 -383 -770 -349
rect 770 -383 866 -349
<< viali >>
rect -605 247 -571 281
rect -409 247 -375 281
rect -213 247 -179 281
rect -17 247 17 281
rect 179 247 213 281
rect 375 247 409 281
rect 571 247 605 281
rect -752 -188 -718 188
rect -654 -188 -620 188
rect -556 -188 -522 188
rect -458 -188 -424 188
rect -360 -188 -326 188
rect -262 -188 -228 188
rect -164 -188 -130 188
rect -66 -188 -32 188
rect 32 -188 66 188
rect 130 -188 164 188
rect 228 -188 262 188
rect 326 -188 360 188
rect 424 -188 458 188
rect 522 -188 556 188
rect 620 -188 654 188
rect 718 -188 752 188
rect -703 -281 -669 -247
rect -507 -281 -473 -247
rect -311 -281 -277 -247
rect -115 -281 -81 -247
rect 81 -281 115 -247
rect 277 -281 311 -247
rect 473 -281 507 -247
rect 669 -281 703 -247
<< metal1 >>
rect -617 281 -559 287
rect -617 247 -605 281
rect -571 247 -559 281
rect -617 241 -559 247
rect -421 281 -363 287
rect -421 247 -409 281
rect -375 247 -363 281
rect -421 241 -363 247
rect -225 281 -167 287
rect -225 247 -213 281
rect -179 247 -167 281
rect -225 241 -167 247
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect 167 281 225 287
rect 167 247 179 281
rect 213 247 225 281
rect 167 241 225 247
rect 363 281 421 287
rect 363 247 375 281
rect 409 247 421 281
rect 363 241 421 247
rect 559 281 617 287
rect 559 247 571 281
rect 605 247 617 281
rect 559 241 617 247
rect -758 188 -712 200
rect -758 -188 -752 188
rect -718 -188 -712 188
rect -758 -200 -712 -188
rect -660 188 -614 200
rect -660 -188 -654 188
rect -620 -188 -614 188
rect -660 -200 -614 -188
rect -562 188 -516 200
rect -562 -188 -556 188
rect -522 -188 -516 188
rect -562 -200 -516 -188
rect -464 188 -418 200
rect -464 -188 -458 188
rect -424 -188 -418 188
rect -464 -200 -418 -188
rect -366 188 -320 200
rect -366 -188 -360 188
rect -326 -188 -320 188
rect -366 -200 -320 -188
rect -268 188 -222 200
rect -268 -188 -262 188
rect -228 -188 -222 188
rect -268 -200 -222 -188
rect -170 188 -124 200
rect -170 -188 -164 188
rect -130 -188 -124 188
rect -170 -200 -124 -188
rect -72 188 -26 200
rect -72 -188 -66 188
rect -32 -188 -26 188
rect -72 -200 -26 -188
rect 26 188 72 200
rect 26 -188 32 188
rect 66 -188 72 188
rect 26 -200 72 -188
rect 124 188 170 200
rect 124 -188 130 188
rect 164 -188 170 188
rect 124 -200 170 -188
rect 222 188 268 200
rect 222 -188 228 188
rect 262 -188 268 188
rect 222 -200 268 -188
rect 320 188 366 200
rect 320 -188 326 188
rect 360 -188 366 188
rect 320 -200 366 -188
rect 418 188 464 200
rect 418 -188 424 188
rect 458 -188 464 188
rect 418 -200 464 -188
rect 516 188 562 200
rect 516 -188 522 188
rect 556 -188 562 188
rect 516 -200 562 -188
rect 614 188 660 200
rect 614 -188 620 188
rect 654 -188 660 188
rect 614 -200 660 -188
rect 712 188 758 200
rect 712 -188 718 188
rect 752 -188 758 188
rect 712 -200 758 -188
rect -715 -247 -657 -241
rect -715 -281 -703 -247
rect -669 -281 -657 -247
rect -715 -287 -657 -281
rect -519 -247 -461 -241
rect -519 -281 -507 -247
rect -473 -281 -461 -247
rect -519 -287 -461 -281
rect -323 -247 -265 -241
rect -323 -281 -311 -247
rect -277 -281 -265 -247
rect -323 -287 -265 -281
rect -127 -247 -69 -241
rect -127 -281 -115 -247
rect -81 -281 -69 -247
rect -127 -287 -69 -281
rect 69 -247 127 -241
rect 69 -281 81 -247
rect 115 -281 127 -247
rect 69 -287 127 -281
rect 265 -247 323 -241
rect 265 -281 277 -247
rect 311 -281 323 -247
rect 265 -287 323 -281
rect 461 -247 519 -241
rect 461 -281 473 -247
rect 507 -281 519 -247
rect 461 -287 519 -281
rect 657 -247 715 -241
rect 657 -281 669 -247
rect 703 -281 715 -247
rect 657 -287 715 -281
<< properties >>
string FIXED_BBOX -849 -366 849 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.2 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
