magic
tech sky130B
magscale 1 2
timestamp 1654683408
<< error_p >>
rect -1325 917 -1267 923
rect -1133 917 -1075 923
rect -941 917 -883 923
rect -749 917 -691 923
rect -557 917 -499 923
rect -365 917 -307 923
rect -173 917 -115 923
rect 19 917 77 923
rect 211 917 269 923
rect 403 917 461 923
rect 595 917 653 923
rect 787 917 845 923
rect 979 917 1037 923
rect 1171 917 1229 923
rect 1363 917 1421 923
rect -1325 883 -1313 917
rect -1133 883 -1121 917
rect -941 883 -929 917
rect -749 883 -737 917
rect -557 883 -545 917
rect -365 883 -353 917
rect -173 883 -161 917
rect 19 883 31 917
rect 211 883 223 917
rect 403 883 415 917
rect 595 883 607 917
rect 787 883 799 917
rect 979 883 991 917
rect 1171 883 1183 917
rect 1363 883 1375 917
rect -1325 877 -1267 883
rect -1133 877 -1075 883
rect -941 877 -883 883
rect -749 877 -691 883
rect -557 877 -499 883
rect -365 877 -307 883
rect -173 877 -115 883
rect 19 877 77 883
rect 211 877 269 883
rect 403 877 461 883
rect 595 877 653 883
rect 787 877 845 883
rect 979 877 1037 883
rect 1171 877 1229 883
rect 1363 877 1421 883
rect -1421 389 -1363 395
rect -1229 389 -1171 395
rect -1037 389 -979 395
rect -845 389 -787 395
rect -653 389 -595 395
rect -461 389 -403 395
rect -269 389 -211 395
rect -77 389 -19 395
rect 115 389 173 395
rect 307 389 365 395
rect 499 389 557 395
rect 691 389 749 395
rect 883 389 941 395
rect 1075 389 1133 395
rect 1267 389 1325 395
rect -1421 355 -1409 389
rect -1229 355 -1217 389
rect -1037 355 -1025 389
rect -845 355 -833 389
rect -653 355 -641 389
rect -461 355 -449 389
rect -269 355 -257 389
rect -77 355 -65 389
rect 115 355 127 389
rect 307 355 319 389
rect 499 355 511 389
rect 691 355 703 389
rect 883 355 895 389
rect 1075 355 1087 389
rect 1267 355 1279 389
rect -1421 349 -1363 355
rect -1229 349 -1171 355
rect -1037 349 -979 355
rect -845 349 -787 355
rect -653 349 -595 355
rect -461 349 -403 355
rect -269 349 -211 355
rect -77 349 -19 355
rect 115 349 173 355
rect 307 349 365 355
rect 499 349 557 355
rect 691 349 749 355
rect 883 349 941 355
rect 1075 349 1133 355
rect 1267 349 1325 355
rect -1421 281 -1363 287
rect -1229 281 -1171 287
rect -1037 281 -979 287
rect -845 281 -787 287
rect -653 281 -595 287
rect -461 281 -403 287
rect -269 281 -211 287
rect -77 281 -19 287
rect 115 281 173 287
rect 307 281 365 287
rect 499 281 557 287
rect 691 281 749 287
rect 883 281 941 287
rect 1075 281 1133 287
rect 1267 281 1325 287
rect -1421 247 -1409 281
rect -1229 247 -1217 281
rect -1037 247 -1025 281
rect -845 247 -833 281
rect -653 247 -641 281
rect -461 247 -449 281
rect -269 247 -257 281
rect -77 247 -65 281
rect 115 247 127 281
rect 307 247 319 281
rect 499 247 511 281
rect 691 247 703 281
rect 883 247 895 281
rect 1075 247 1087 281
rect 1267 247 1279 281
rect -1421 241 -1363 247
rect -1229 241 -1171 247
rect -1037 241 -979 247
rect -845 241 -787 247
rect -653 241 -595 247
rect -461 241 -403 247
rect -269 241 -211 247
rect -77 241 -19 247
rect 115 241 173 247
rect 307 241 365 247
rect 499 241 557 247
rect 691 241 749 247
rect 883 241 941 247
rect 1075 241 1133 247
rect 1267 241 1325 247
rect -1325 -247 -1267 -241
rect -1133 -247 -1075 -241
rect -941 -247 -883 -241
rect -749 -247 -691 -241
rect -557 -247 -499 -241
rect -365 -247 -307 -241
rect -173 -247 -115 -241
rect 19 -247 77 -241
rect 211 -247 269 -241
rect 403 -247 461 -241
rect 595 -247 653 -241
rect 787 -247 845 -241
rect 979 -247 1037 -241
rect 1171 -247 1229 -241
rect 1363 -247 1421 -241
rect -1325 -281 -1313 -247
rect -1133 -281 -1121 -247
rect -941 -281 -929 -247
rect -749 -281 -737 -247
rect -557 -281 -545 -247
rect -365 -281 -353 -247
rect -173 -281 -161 -247
rect 19 -281 31 -247
rect 211 -281 223 -247
rect 403 -281 415 -247
rect 595 -281 607 -247
rect 787 -281 799 -247
rect 979 -281 991 -247
rect 1171 -281 1183 -247
rect 1363 -281 1375 -247
rect -1325 -287 -1267 -281
rect -1133 -287 -1075 -281
rect -941 -287 -883 -281
rect -749 -287 -691 -281
rect -557 -287 -499 -281
rect -365 -287 -307 -281
rect -173 -287 -115 -281
rect 19 -287 77 -281
rect 211 -287 269 -281
rect 403 -287 461 -281
rect 595 -287 653 -281
rect 787 -287 845 -281
rect 979 -287 1037 -281
rect 1171 -287 1229 -281
rect 1363 -287 1421 -281
rect -1325 -355 -1267 -349
rect -1133 -355 -1075 -349
rect -941 -355 -883 -349
rect -749 -355 -691 -349
rect -557 -355 -499 -349
rect -365 -355 -307 -349
rect -173 -355 -115 -349
rect 19 -355 77 -349
rect 211 -355 269 -349
rect 403 -355 461 -349
rect 595 -355 653 -349
rect 787 -355 845 -349
rect 979 -355 1037 -349
rect 1171 -355 1229 -349
rect 1363 -355 1421 -349
rect -1325 -389 -1313 -355
rect -1133 -389 -1121 -355
rect -941 -389 -929 -355
rect -749 -389 -737 -355
rect -557 -389 -545 -355
rect -365 -389 -353 -355
rect -173 -389 -161 -355
rect 19 -389 31 -355
rect 211 -389 223 -355
rect 403 -389 415 -355
rect 595 -389 607 -355
rect 787 -389 799 -355
rect 979 -389 991 -355
rect 1171 -389 1183 -355
rect 1363 -389 1375 -355
rect -1325 -395 -1267 -389
rect -1133 -395 -1075 -389
rect -941 -395 -883 -389
rect -749 -395 -691 -389
rect -557 -395 -499 -389
rect -365 -395 -307 -389
rect -173 -395 -115 -389
rect 19 -395 77 -389
rect 211 -395 269 -389
rect 403 -395 461 -389
rect 595 -395 653 -389
rect 787 -395 845 -389
rect 979 -395 1037 -389
rect 1171 -395 1229 -389
rect 1363 -395 1421 -389
rect -1421 -883 -1363 -877
rect -1229 -883 -1171 -877
rect -1037 -883 -979 -877
rect -845 -883 -787 -877
rect -653 -883 -595 -877
rect -461 -883 -403 -877
rect -269 -883 -211 -877
rect -77 -883 -19 -877
rect 115 -883 173 -877
rect 307 -883 365 -877
rect 499 -883 557 -877
rect 691 -883 749 -877
rect 883 -883 941 -877
rect 1075 -883 1133 -877
rect 1267 -883 1325 -877
rect -1421 -917 -1409 -883
rect -1229 -917 -1217 -883
rect -1037 -917 -1025 -883
rect -845 -917 -833 -883
rect -653 -917 -641 -883
rect -461 -917 -449 -883
rect -269 -917 -257 -883
rect -77 -917 -65 -883
rect 115 -917 127 -883
rect 307 -917 319 -883
rect 499 -917 511 -883
rect 691 -917 703 -883
rect 883 -917 895 -883
rect 1075 -917 1087 -883
rect 1267 -917 1279 -883
rect -1421 -923 -1363 -917
rect -1229 -923 -1171 -917
rect -1037 -923 -979 -917
rect -845 -923 -787 -917
rect -653 -923 -595 -917
rect -461 -923 -403 -917
rect -269 -923 -211 -917
rect -77 -923 -19 -917
rect 115 -923 173 -917
rect 307 -923 365 -917
rect 499 -923 557 -917
rect 691 -923 749 -917
rect 883 -923 941 -917
rect 1075 -923 1133 -917
rect 1267 -923 1325 -917
<< nwell >>
rect -1607 -1055 1607 1055
<< pmos >>
rect -1407 436 -1377 836
rect -1311 436 -1281 836
rect -1215 436 -1185 836
rect -1119 436 -1089 836
rect -1023 436 -993 836
rect -927 436 -897 836
rect -831 436 -801 836
rect -735 436 -705 836
rect -639 436 -609 836
rect -543 436 -513 836
rect -447 436 -417 836
rect -351 436 -321 836
rect -255 436 -225 836
rect -159 436 -129 836
rect -63 436 -33 836
rect 33 436 63 836
rect 129 436 159 836
rect 225 436 255 836
rect 321 436 351 836
rect 417 436 447 836
rect 513 436 543 836
rect 609 436 639 836
rect 705 436 735 836
rect 801 436 831 836
rect 897 436 927 836
rect 993 436 1023 836
rect 1089 436 1119 836
rect 1185 436 1215 836
rect 1281 436 1311 836
rect 1377 436 1407 836
rect -1407 -200 -1377 200
rect -1311 -200 -1281 200
rect -1215 -200 -1185 200
rect -1119 -200 -1089 200
rect -1023 -200 -993 200
rect -927 -200 -897 200
rect -831 -200 -801 200
rect -735 -200 -705 200
rect -639 -200 -609 200
rect -543 -200 -513 200
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect 513 -200 543 200
rect 609 -200 639 200
rect 705 -200 735 200
rect 801 -200 831 200
rect 897 -200 927 200
rect 993 -200 1023 200
rect 1089 -200 1119 200
rect 1185 -200 1215 200
rect 1281 -200 1311 200
rect 1377 -200 1407 200
rect -1407 -836 -1377 -436
rect -1311 -836 -1281 -436
rect -1215 -836 -1185 -436
rect -1119 -836 -1089 -436
rect -1023 -836 -993 -436
rect -927 -836 -897 -436
rect -831 -836 -801 -436
rect -735 -836 -705 -436
rect -639 -836 -609 -436
rect -543 -836 -513 -436
rect -447 -836 -417 -436
rect -351 -836 -321 -436
rect -255 -836 -225 -436
rect -159 -836 -129 -436
rect -63 -836 -33 -436
rect 33 -836 63 -436
rect 129 -836 159 -436
rect 225 -836 255 -436
rect 321 -836 351 -436
rect 417 -836 447 -436
rect 513 -836 543 -436
rect 609 -836 639 -436
rect 705 -836 735 -436
rect 801 -836 831 -436
rect 897 -836 927 -436
rect 993 -836 1023 -436
rect 1089 -836 1119 -436
rect 1185 -836 1215 -436
rect 1281 -836 1311 -436
rect 1377 -836 1407 -436
<< pdiff >>
rect -1469 824 -1407 836
rect -1469 448 -1457 824
rect -1423 448 -1407 824
rect -1469 436 -1407 448
rect -1377 824 -1311 836
rect -1377 448 -1361 824
rect -1327 448 -1311 824
rect -1377 436 -1311 448
rect -1281 824 -1215 836
rect -1281 448 -1265 824
rect -1231 448 -1215 824
rect -1281 436 -1215 448
rect -1185 824 -1119 836
rect -1185 448 -1169 824
rect -1135 448 -1119 824
rect -1185 436 -1119 448
rect -1089 824 -1023 836
rect -1089 448 -1073 824
rect -1039 448 -1023 824
rect -1089 436 -1023 448
rect -993 824 -927 836
rect -993 448 -977 824
rect -943 448 -927 824
rect -993 436 -927 448
rect -897 824 -831 836
rect -897 448 -881 824
rect -847 448 -831 824
rect -897 436 -831 448
rect -801 824 -735 836
rect -801 448 -785 824
rect -751 448 -735 824
rect -801 436 -735 448
rect -705 824 -639 836
rect -705 448 -689 824
rect -655 448 -639 824
rect -705 436 -639 448
rect -609 824 -543 836
rect -609 448 -593 824
rect -559 448 -543 824
rect -609 436 -543 448
rect -513 824 -447 836
rect -513 448 -497 824
rect -463 448 -447 824
rect -513 436 -447 448
rect -417 824 -351 836
rect -417 448 -401 824
rect -367 448 -351 824
rect -417 436 -351 448
rect -321 824 -255 836
rect -321 448 -305 824
rect -271 448 -255 824
rect -321 436 -255 448
rect -225 824 -159 836
rect -225 448 -209 824
rect -175 448 -159 824
rect -225 436 -159 448
rect -129 824 -63 836
rect -129 448 -113 824
rect -79 448 -63 824
rect -129 436 -63 448
rect -33 824 33 836
rect -33 448 -17 824
rect 17 448 33 824
rect -33 436 33 448
rect 63 824 129 836
rect 63 448 79 824
rect 113 448 129 824
rect 63 436 129 448
rect 159 824 225 836
rect 159 448 175 824
rect 209 448 225 824
rect 159 436 225 448
rect 255 824 321 836
rect 255 448 271 824
rect 305 448 321 824
rect 255 436 321 448
rect 351 824 417 836
rect 351 448 367 824
rect 401 448 417 824
rect 351 436 417 448
rect 447 824 513 836
rect 447 448 463 824
rect 497 448 513 824
rect 447 436 513 448
rect 543 824 609 836
rect 543 448 559 824
rect 593 448 609 824
rect 543 436 609 448
rect 639 824 705 836
rect 639 448 655 824
rect 689 448 705 824
rect 639 436 705 448
rect 735 824 801 836
rect 735 448 751 824
rect 785 448 801 824
rect 735 436 801 448
rect 831 824 897 836
rect 831 448 847 824
rect 881 448 897 824
rect 831 436 897 448
rect 927 824 993 836
rect 927 448 943 824
rect 977 448 993 824
rect 927 436 993 448
rect 1023 824 1089 836
rect 1023 448 1039 824
rect 1073 448 1089 824
rect 1023 436 1089 448
rect 1119 824 1185 836
rect 1119 448 1135 824
rect 1169 448 1185 824
rect 1119 436 1185 448
rect 1215 824 1281 836
rect 1215 448 1231 824
rect 1265 448 1281 824
rect 1215 436 1281 448
rect 1311 824 1377 836
rect 1311 448 1327 824
rect 1361 448 1377 824
rect 1311 436 1377 448
rect 1407 824 1469 836
rect 1407 448 1423 824
rect 1457 448 1469 824
rect 1407 436 1469 448
rect -1469 188 -1407 200
rect -1469 -188 -1457 188
rect -1423 -188 -1407 188
rect -1469 -200 -1407 -188
rect -1377 188 -1311 200
rect -1377 -188 -1361 188
rect -1327 -188 -1311 188
rect -1377 -200 -1311 -188
rect -1281 188 -1215 200
rect -1281 -188 -1265 188
rect -1231 -188 -1215 188
rect -1281 -200 -1215 -188
rect -1185 188 -1119 200
rect -1185 -188 -1169 188
rect -1135 -188 -1119 188
rect -1185 -200 -1119 -188
rect -1089 188 -1023 200
rect -1089 -188 -1073 188
rect -1039 -188 -1023 188
rect -1089 -200 -1023 -188
rect -993 188 -927 200
rect -993 -188 -977 188
rect -943 -188 -927 188
rect -993 -200 -927 -188
rect -897 188 -831 200
rect -897 -188 -881 188
rect -847 -188 -831 188
rect -897 -200 -831 -188
rect -801 188 -735 200
rect -801 -188 -785 188
rect -751 -188 -735 188
rect -801 -200 -735 -188
rect -705 188 -639 200
rect -705 -188 -689 188
rect -655 -188 -639 188
rect -705 -200 -639 -188
rect -609 188 -543 200
rect -609 -188 -593 188
rect -559 -188 -543 188
rect -609 -200 -543 -188
rect -513 188 -447 200
rect -513 -188 -497 188
rect -463 -188 -447 188
rect -513 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 513 200
rect 447 -188 463 188
rect 497 -188 513 188
rect 447 -200 513 -188
rect 543 188 609 200
rect 543 -188 559 188
rect 593 -188 609 188
rect 543 -200 609 -188
rect 639 188 705 200
rect 639 -188 655 188
rect 689 -188 705 188
rect 639 -200 705 -188
rect 735 188 801 200
rect 735 -188 751 188
rect 785 -188 801 188
rect 735 -200 801 -188
rect 831 188 897 200
rect 831 -188 847 188
rect 881 -188 897 188
rect 831 -200 897 -188
rect 927 188 993 200
rect 927 -188 943 188
rect 977 -188 993 188
rect 927 -200 993 -188
rect 1023 188 1089 200
rect 1023 -188 1039 188
rect 1073 -188 1089 188
rect 1023 -200 1089 -188
rect 1119 188 1185 200
rect 1119 -188 1135 188
rect 1169 -188 1185 188
rect 1119 -200 1185 -188
rect 1215 188 1281 200
rect 1215 -188 1231 188
rect 1265 -188 1281 188
rect 1215 -200 1281 -188
rect 1311 188 1377 200
rect 1311 -188 1327 188
rect 1361 -188 1377 188
rect 1311 -200 1377 -188
rect 1407 188 1469 200
rect 1407 -188 1423 188
rect 1457 -188 1469 188
rect 1407 -200 1469 -188
rect -1469 -448 -1407 -436
rect -1469 -824 -1457 -448
rect -1423 -824 -1407 -448
rect -1469 -836 -1407 -824
rect -1377 -448 -1311 -436
rect -1377 -824 -1361 -448
rect -1327 -824 -1311 -448
rect -1377 -836 -1311 -824
rect -1281 -448 -1215 -436
rect -1281 -824 -1265 -448
rect -1231 -824 -1215 -448
rect -1281 -836 -1215 -824
rect -1185 -448 -1119 -436
rect -1185 -824 -1169 -448
rect -1135 -824 -1119 -448
rect -1185 -836 -1119 -824
rect -1089 -448 -1023 -436
rect -1089 -824 -1073 -448
rect -1039 -824 -1023 -448
rect -1089 -836 -1023 -824
rect -993 -448 -927 -436
rect -993 -824 -977 -448
rect -943 -824 -927 -448
rect -993 -836 -927 -824
rect -897 -448 -831 -436
rect -897 -824 -881 -448
rect -847 -824 -831 -448
rect -897 -836 -831 -824
rect -801 -448 -735 -436
rect -801 -824 -785 -448
rect -751 -824 -735 -448
rect -801 -836 -735 -824
rect -705 -448 -639 -436
rect -705 -824 -689 -448
rect -655 -824 -639 -448
rect -705 -836 -639 -824
rect -609 -448 -543 -436
rect -609 -824 -593 -448
rect -559 -824 -543 -448
rect -609 -836 -543 -824
rect -513 -448 -447 -436
rect -513 -824 -497 -448
rect -463 -824 -447 -448
rect -513 -836 -447 -824
rect -417 -448 -351 -436
rect -417 -824 -401 -448
rect -367 -824 -351 -448
rect -417 -836 -351 -824
rect -321 -448 -255 -436
rect -321 -824 -305 -448
rect -271 -824 -255 -448
rect -321 -836 -255 -824
rect -225 -448 -159 -436
rect -225 -824 -209 -448
rect -175 -824 -159 -448
rect -225 -836 -159 -824
rect -129 -448 -63 -436
rect -129 -824 -113 -448
rect -79 -824 -63 -448
rect -129 -836 -63 -824
rect -33 -448 33 -436
rect -33 -824 -17 -448
rect 17 -824 33 -448
rect -33 -836 33 -824
rect 63 -448 129 -436
rect 63 -824 79 -448
rect 113 -824 129 -448
rect 63 -836 129 -824
rect 159 -448 225 -436
rect 159 -824 175 -448
rect 209 -824 225 -448
rect 159 -836 225 -824
rect 255 -448 321 -436
rect 255 -824 271 -448
rect 305 -824 321 -448
rect 255 -836 321 -824
rect 351 -448 417 -436
rect 351 -824 367 -448
rect 401 -824 417 -448
rect 351 -836 417 -824
rect 447 -448 513 -436
rect 447 -824 463 -448
rect 497 -824 513 -448
rect 447 -836 513 -824
rect 543 -448 609 -436
rect 543 -824 559 -448
rect 593 -824 609 -448
rect 543 -836 609 -824
rect 639 -448 705 -436
rect 639 -824 655 -448
rect 689 -824 705 -448
rect 639 -836 705 -824
rect 735 -448 801 -436
rect 735 -824 751 -448
rect 785 -824 801 -448
rect 735 -836 801 -824
rect 831 -448 897 -436
rect 831 -824 847 -448
rect 881 -824 897 -448
rect 831 -836 897 -824
rect 927 -448 993 -436
rect 927 -824 943 -448
rect 977 -824 993 -448
rect 927 -836 993 -824
rect 1023 -448 1089 -436
rect 1023 -824 1039 -448
rect 1073 -824 1089 -448
rect 1023 -836 1089 -824
rect 1119 -448 1185 -436
rect 1119 -824 1135 -448
rect 1169 -824 1185 -448
rect 1119 -836 1185 -824
rect 1215 -448 1281 -436
rect 1215 -824 1231 -448
rect 1265 -824 1281 -448
rect 1215 -836 1281 -824
rect 1311 -448 1377 -436
rect 1311 -824 1327 -448
rect 1361 -824 1377 -448
rect 1311 -836 1377 -824
rect 1407 -448 1469 -436
rect 1407 -824 1423 -448
rect 1457 -824 1469 -448
rect 1407 -836 1469 -824
<< pdiffc >>
rect -1457 448 -1423 824
rect -1361 448 -1327 824
rect -1265 448 -1231 824
rect -1169 448 -1135 824
rect -1073 448 -1039 824
rect -977 448 -943 824
rect -881 448 -847 824
rect -785 448 -751 824
rect -689 448 -655 824
rect -593 448 -559 824
rect -497 448 -463 824
rect -401 448 -367 824
rect -305 448 -271 824
rect -209 448 -175 824
rect -113 448 -79 824
rect -17 448 17 824
rect 79 448 113 824
rect 175 448 209 824
rect 271 448 305 824
rect 367 448 401 824
rect 463 448 497 824
rect 559 448 593 824
rect 655 448 689 824
rect 751 448 785 824
rect 847 448 881 824
rect 943 448 977 824
rect 1039 448 1073 824
rect 1135 448 1169 824
rect 1231 448 1265 824
rect 1327 448 1361 824
rect 1423 448 1457 824
rect -1457 -188 -1423 188
rect -1361 -188 -1327 188
rect -1265 -188 -1231 188
rect -1169 -188 -1135 188
rect -1073 -188 -1039 188
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect 1039 -188 1073 188
rect 1135 -188 1169 188
rect 1231 -188 1265 188
rect 1327 -188 1361 188
rect 1423 -188 1457 188
rect -1457 -824 -1423 -448
rect -1361 -824 -1327 -448
rect -1265 -824 -1231 -448
rect -1169 -824 -1135 -448
rect -1073 -824 -1039 -448
rect -977 -824 -943 -448
rect -881 -824 -847 -448
rect -785 -824 -751 -448
rect -689 -824 -655 -448
rect -593 -824 -559 -448
rect -497 -824 -463 -448
rect -401 -824 -367 -448
rect -305 -824 -271 -448
rect -209 -824 -175 -448
rect -113 -824 -79 -448
rect -17 -824 17 -448
rect 79 -824 113 -448
rect 175 -824 209 -448
rect 271 -824 305 -448
rect 367 -824 401 -448
rect 463 -824 497 -448
rect 559 -824 593 -448
rect 655 -824 689 -448
rect 751 -824 785 -448
rect 847 -824 881 -448
rect 943 -824 977 -448
rect 1039 -824 1073 -448
rect 1135 -824 1169 -448
rect 1231 -824 1265 -448
rect 1327 -824 1361 -448
rect 1423 -824 1457 -448
<< nsubdiff >>
rect -1571 985 -1475 1019
rect 1475 985 1571 1019
rect -1571 923 -1537 985
rect 1537 923 1571 985
rect -1571 -985 -1537 -923
rect 1537 -985 1571 -923
rect -1571 -1019 -1475 -985
rect 1475 -1019 1571 -985
<< nsubdiffcont >>
rect -1475 985 1475 1019
rect -1571 -923 -1537 923
rect 1537 -923 1571 923
rect -1475 -1019 1475 -985
<< poly >>
rect -1329 917 -1263 933
rect -1329 883 -1313 917
rect -1279 883 -1263 917
rect -1329 867 -1263 883
rect -1137 917 -1071 933
rect -1137 883 -1121 917
rect -1087 883 -1071 917
rect -1137 867 -1071 883
rect -945 917 -879 933
rect -945 883 -929 917
rect -895 883 -879 917
rect -945 867 -879 883
rect -753 917 -687 933
rect -753 883 -737 917
rect -703 883 -687 917
rect -753 867 -687 883
rect -561 917 -495 933
rect -561 883 -545 917
rect -511 883 -495 917
rect -561 867 -495 883
rect -369 917 -303 933
rect -369 883 -353 917
rect -319 883 -303 917
rect -369 867 -303 883
rect -177 917 -111 933
rect -177 883 -161 917
rect -127 883 -111 917
rect -177 867 -111 883
rect 15 917 81 933
rect 15 883 31 917
rect 65 883 81 917
rect 15 867 81 883
rect 207 917 273 933
rect 207 883 223 917
rect 257 883 273 917
rect 207 867 273 883
rect 399 917 465 933
rect 399 883 415 917
rect 449 883 465 917
rect 399 867 465 883
rect 591 917 657 933
rect 591 883 607 917
rect 641 883 657 917
rect 591 867 657 883
rect 783 917 849 933
rect 783 883 799 917
rect 833 883 849 917
rect 783 867 849 883
rect 975 917 1041 933
rect 975 883 991 917
rect 1025 883 1041 917
rect 975 867 1041 883
rect 1167 917 1233 933
rect 1167 883 1183 917
rect 1217 883 1233 917
rect 1167 867 1233 883
rect 1359 917 1425 933
rect 1359 883 1375 917
rect 1409 883 1425 917
rect 1359 867 1425 883
rect -1407 836 -1377 862
rect -1311 836 -1281 867
rect -1215 836 -1185 862
rect -1119 836 -1089 867
rect -1023 836 -993 862
rect -927 836 -897 867
rect -831 836 -801 862
rect -735 836 -705 867
rect -639 836 -609 862
rect -543 836 -513 867
rect -447 836 -417 862
rect -351 836 -321 867
rect -255 836 -225 862
rect -159 836 -129 867
rect -63 836 -33 862
rect 33 836 63 867
rect 129 836 159 862
rect 225 836 255 867
rect 321 836 351 862
rect 417 836 447 867
rect 513 836 543 862
rect 609 836 639 867
rect 705 836 735 862
rect 801 836 831 867
rect 897 836 927 862
rect 993 836 1023 867
rect 1089 836 1119 862
rect 1185 836 1215 867
rect 1281 836 1311 862
rect 1377 836 1407 867
rect -1407 405 -1377 436
rect -1311 410 -1281 436
rect -1215 405 -1185 436
rect -1119 410 -1089 436
rect -1023 405 -993 436
rect -927 410 -897 436
rect -831 405 -801 436
rect -735 410 -705 436
rect -639 405 -609 436
rect -543 410 -513 436
rect -447 405 -417 436
rect -351 410 -321 436
rect -255 405 -225 436
rect -159 410 -129 436
rect -63 405 -33 436
rect 33 410 63 436
rect 129 405 159 436
rect 225 410 255 436
rect 321 405 351 436
rect 417 410 447 436
rect 513 405 543 436
rect 609 410 639 436
rect 705 405 735 436
rect 801 410 831 436
rect 897 405 927 436
rect 993 410 1023 436
rect 1089 405 1119 436
rect 1185 410 1215 436
rect 1281 405 1311 436
rect 1377 410 1407 436
rect -1425 389 -1359 405
rect -1425 355 -1409 389
rect -1375 355 -1359 389
rect -1425 339 -1359 355
rect -1233 389 -1167 405
rect -1233 355 -1217 389
rect -1183 355 -1167 389
rect -1233 339 -1167 355
rect -1041 389 -975 405
rect -1041 355 -1025 389
rect -991 355 -975 389
rect -1041 339 -975 355
rect -849 389 -783 405
rect -849 355 -833 389
rect -799 355 -783 389
rect -849 339 -783 355
rect -657 389 -591 405
rect -657 355 -641 389
rect -607 355 -591 389
rect -657 339 -591 355
rect -465 389 -399 405
rect -465 355 -449 389
rect -415 355 -399 389
rect -465 339 -399 355
rect -273 389 -207 405
rect -273 355 -257 389
rect -223 355 -207 389
rect -273 339 -207 355
rect -81 389 -15 405
rect -81 355 -65 389
rect -31 355 -15 389
rect -81 339 -15 355
rect 111 389 177 405
rect 111 355 127 389
rect 161 355 177 389
rect 111 339 177 355
rect 303 389 369 405
rect 303 355 319 389
rect 353 355 369 389
rect 303 339 369 355
rect 495 389 561 405
rect 495 355 511 389
rect 545 355 561 389
rect 495 339 561 355
rect 687 389 753 405
rect 687 355 703 389
rect 737 355 753 389
rect 687 339 753 355
rect 879 389 945 405
rect 879 355 895 389
rect 929 355 945 389
rect 879 339 945 355
rect 1071 389 1137 405
rect 1071 355 1087 389
rect 1121 355 1137 389
rect 1071 339 1137 355
rect 1263 389 1329 405
rect 1263 355 1279 389
rect 1313 355 1329 389
rect 1263 339 1329 355
rect -1425 281 -1359 297
rect -1425 247 -1409 281
rect -1375 247 -1359 281
rect -1425 231 -1359 247
rect -1233 281 -1167 297
rect -1233 247 -1217 281
rect -1183 247 -1167 281
rect -1233 231 -1167 247
rect -1041 281 -975 297
rect -1041 247 -1025 281
rect -991 247 -975 281
rect -1041 231 -975 247
rect -849 281 -783 297
rect -849 247 -833 281
rect -799 247 -783 281
rect -849 231 -783 247
rect -657 281 -591 297
rect -657 247 -641 281
rect -607 247 -591 281
rect -657 231 -591 247
rect -465 281 -399 297
rect -465 247 -449 281
rect -415 247 -399 281
rect -465 231 -399 247
rect -273 281 -207 297
rect -273 247 -257 281
rect -223 247 -207 281
rect -273 231 -207 247
rect -81 281 -15 297
rect -81 247 -65 281
rect -31 247 -15 281
rect -81 231 -15 247
rect 111 281 177 297
rect 111 247 127 281
rect 161 247 177 281
rect 111 231 177 247
rect 303 281 369 297
rect 303 247 319 281
rect 353 247 369 281
rect 303 231 369 247
rect 495 281 561 297
rect 495 247 511 281
rect 545 247 561 281
rect 495 231 561 247
rect 687 281 753 297
rect 687 247 703 281
rect 737 247 753 281
rect 687 231 753 247
rect 879 281 945 297
rect 879 247 895 281
rect 929 247 945 281
rect 879 231 945 247
rect 1071 281 1137 297
rect 1071 247 1087 281
rect 1121 247 1137 281
rect 1071 231 1137 247
rect 1263 281 1329 297
rect 1263 247 1279 281
rect 1313 247 1329 281
rect 1263 231 1329 247
rect -1407 200 -1377 231
rect -1311 200 -1281 226
rect -1215 200 -1185 231
rect -1119 200 -1089 226
rect -1023 200 -993 231
rect -927 200 -897 226
rect -831 200 -801 231
rect -735 200 -705 226
rect -639 200 -609 231
rect -543 200 -513 226
rect -447 200 -417 231
rect -351 200 -321 226
rect -255 200 -225 231
rect -159 200 -129 226
rect -63 200 -33 231
rect 33 200 63 226
rect 129 200 159 231
rect 225 200 255 226
rect 321 200 351 231
rect 417 200 447 226
rect 513 200 543 231
rect 609 200 639 226
rect 705 200 735 231
rect 801 200 831 226
rect 897 200 927 231
rect 993 200 1023 226
rect 1089 200 1119 231
rect 1185 200 1215 226
rect 1281 200 1311 231
rect 1377 200 1407 226
rect -1407 -226 -1377 -200
rect -1311 -231 -1281 -200
rect -1215 -226 -1185 -200
rect -1119 -231 -1089 -200
rect -1023 -226 -993 -200
rect -927 -231 -897 -200
rect -831 -226 -801 -200
rect -735 -231 -705 -200
rect -639 -226 -609 -200
rect -543 -231 -513 -200
rect -447 -226 -417 -200
rect -351 -231 -321 -200
rect -255 -226 -225 -200
rect -159 -231 -129 -200
rect -63 -226 -33 -200
rect 33 -231 63 -200
rect 129 -226 159 -200
rect 225 -231 255 -200
rect 321 -226 351 -200
rect 417 -231 447 -200
rect 513 -226 543 -200
rect 609 -231 639 -200
rect 705 -226 735 -200
rect 801 -231 831 -200
rect 897 -226 927 -200
rect 993 -231 1023 -200
rect 1089 -226 1119 -200
rect 1185 -231 1215 -200
rect 1281 -226 1311 -200
rect 1377 -231 1407 -200
rect -1329 -247 -1263 -231
rect -1329 -281 -1313 -247
rect -1279 -281 -1263 -247
rect -1329 -297 -1263 -281
rect -1137 -247 -1071 -231
rect -1137 -281 -1121 -247
rect -1087 -281 -1071 -247
rect -1137 -297 -1071 -281
rect -945 -247 -879 -231
rect -945 -281 -929 -247
rect -895 -281 -879 -247
rect -945 -297 -879 -281
rect -753 -247 -687 -231
rect -753 -281 -737 -247
rect -703 -281 -687 -247
rect -753 -297 -687 -281
rect -561 -247 -495 -231
rect -561 -281 -545 -247
rect -511 -281 -495 -247
rect -561 -297 -495 -281
rect -369 -247 -303 -231
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -369 -297 -303 -281
rect -177 -247 -111 -231
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect -177 -297 -111 -281
rect 15 -247 81 -231
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 15 -297 81 -281
rect 207 -247 273 -231
rect 207 -281 223 -247
rect 257 -281 273 -247
rect 207 -297 273 -281
rect 399 -247 465 -231
rect 399 -281 415 -247
rect 449 -281 465 -247
rect 399 -297 465 -281
rect 591 -247 657 -231
rect 591 -281 607 -247
rect 641 -281 657 -247
rect 591 -297 657 -281
rect 783 -247 849 -231
rect 783 -281 799 -247
rect 833 -281 849 -247
rect 783 -297 849 -281
rect 975 -247 1041 -231
rect 975 -281 991 -247
rect 1025 -281 1041 -247
rect 975 -297 1041 -281
rect 1167 -247 1233 -231
rect 1167 -281 1183 -247
rect 1217 -281 1233 -247
rect 1167 -297 1233 -281
rect 1359 -247 1425 -231
rect 1359 -281 1375 -247
rect 1409 -281 1425 -247
rect 1359 -297 1425 -281
rect -1329 -355 -1263 -339
rect -1329 -389 -1313 -355
rect -1279 -389 -1263 -355
rect -1329 -405 -1263 -389
rect -1137 -355 -1071 -339
rect -1137 -389 -1121 -355
rect -1087 -389 -1071 -355
rect -1137 -405 -1071 -389
rect -945 -355 -879 -339
rect -945 -389 -929 -355
rect -895 -389 -879 -355
rect -945 -405 -879 -389
rect -753 -355 -687 -339
rect -753 -389 -737 -355
rect -703 -389 -687 -355
rect -753 -405 -687 -389
rect -561 -355 -495 -339
rect -561 -389 -545 -355
rect -511 -389 -495 -355
rect -561 -405 -495 -389
rect -369 -355 -303 -339
rect -369 -389 -353 -355
rect -319 -389 -303 -355
rect -369 -405 -303 -389
rect -177 -355 -111 -339
rect -177 -389 -161 -355
rect -127 -389 -111 -355
rect -177 -405 -111 -389
rect 15 -355 81 -339
rect 15 -389 31 -355
rect 65 -389 81 -355
rect 15 -405 81 -389
rect 207 -355 273 -339
rect 207 -389 223 -355
rect 257 -389 273 -355
rect 207 -405 273 -389
rect 399 -355 465 -339
rect 399 -389 415 -355
rect 449 -389 465 -355
rect 399 -405 465 -389
rect 591 -355 657 -339
rect 591 -389 607 -355
rect 641 -389 657 -355
rect 591 -405 657 -389
rect 783 -355 849 -339
rect 783 -389 799 -355
rect 833 -389 849 -355
rect 783 -405 849 -389
rect 975 -355 1041 -339
rect 975 -389 991 -355
rect 1025 -389 1041 -355
rect 975 -405 1041 -389
rect 1167 -355 1233 -339
rect 1167 -389 1183 -355
rect 1217 -389 1233 -355
rect 1167 -405 1233 -389
rect 1359 -355 1425 -339
rect 1359 -389 1375 -355
rect 1409 -389 1425 -355
rect 1359 -405 1425 -389
rect -1407 -436 -1377 -410
rect -1311 -436 -1281 -405
rect -1215 -436 -1185 -410
rect -1119 -436 -1089 -405
rect -1023 -436 -993 -410
rect -927 -436 -897 -405
rect -831 -436 -801 -410
rect -735 -436 -705 -405
rect -639 -436 -609 -410
rect -543 -436 -513 -405
rect -447 -436 -417 -410
rect -351 -436 -321 -405
rect -255 -436 -225 -410
rect -159 -436 -129 -405
rect -63 -436 -33 -410
rect 33 -436 63 -405
rect 129 -436 159 -410
rect 225 -436 255 -405
rect 321 -436 351 -410
rect 417 -436 447 -405
rect 513 -436 543 -410
rect 609 -436 639 -405
rect 705 -436 735 -410
rect 801 -436 831 -405
rect 897 -436 927 -410
rect 993 -436 1023 -405
rect 1089 -436 1119 -410
rect 1185 -436 1215 -405
rect 1281 -436 1311 -410
rect 1377 -436 1407 -405
rect -1407 -867 -1377 -836
rect -1311 -862 -1281 -836
rect -1215 -867 -1185 -836
rect -1119 -862 -1089 -836
rect -1023 -867 -993 -836
rect -927 -862 -897 -836
rect -831 -867 -801 -836
rect -735 -862 -705 -836
rect -639 -867 -609 -836
rect -543 -862 -513 -836
rect -447 -867 -417 -836
rect -351 -862 -321 -836
rect -255 -867 -225 -836
rect -159 -862 -129 -836
rect -63 -867 -33 -836
rect 33 -862 63 -836
rect 129 -867 159 -836
rect 225 -862 255 -836
rect 321 -867 351 -836
rect 417 -862 447 -836
rect 513 -867 543 -836
rect 609 -862 639 -836
rect 705 -867 735 -836
rect 801 -862 831 -836
rect 897 -867 927 -836
rect 993 -862 1023 -836
rect 1089 -867 1119 -836
rect 1185 -862 1215 -836
rect 1281 -867 1311 -836
rect 1377 -862 1407 -836
rect -1425 -883 -1359 -867
rect -1425 -917 -1409 -883
rect -1375 -917 -1359 -883
rect -1425 -933 -1359 -917
rect -1233 -883 -1167 -867
rect -1233 -917 -1217 -883
rect -1183 -917 -1167 -883
rect -1233 -933 -1167 -917
rect -1041 -883 -975 -867
rect -1041 -917 -1025 -883
rect -991 -917 -975 -883
rect -1041 -933 -975 -917
rect -849 -883 -783 -867
rect -849 -917 -833 -883
rect -799 -917 -783 -883
rect -849 -933 -783 -917
rect -657 -883 -591 -867
rect -657 -917 -641 -883
rect -607 -917 -591 -883
rect -657 -933 -591 -917
rect -465 -883 -399 -867
rect -465 -917 -449 -883
rect -415 -917 -399 -883
rect -465 -933 -399 -917
rect -273 -883 -207 -867
rect -273 -917 -257 -883
rect -223 -917 -207 -883
rect -273 -933 -207 -917
rect -81 -883 -15 -867
rect -81 -917 -65 -883
rect -31 -917 -15 -883
rect -81 -933 -15 -917
rect 111 -883 177 -867
rect 111 -917 127 -883
rect 161 -917 177 -883
rect 111 -933 177 -917
rect 303 -883 369 -867
rect 303 -917 319 -883
rect 353 -917 369 -883
rect 303 -933 369 -917
rect 495 -883 561 -867
rect 495 -917 511 -883
rect 545 -917 561 -883
rect 495 -933 561 -917
rect 687 -883 753 -867
rect 687 -917 703 -883
rect 737 -917 753 -883
rect 687 -933 753 -917
rect 879 -883 945 -867
rect 879 -917 895 -883
rect 929 -917 945 -883
rect 879 -933 945 -917
rect 1071 -883 1137 -867
rect 1071 -917 1087 -883
rect 1121 -917 1137 -883
rect 1071 -933 1137 -917
rect 1263 -883 1329 -867
rect 1263 -917 1279 -883
rect 1313 -917 1329 -883
rect 1263 -933 1329 -917
<< polycont >>
rect -1313 883 -1279 917
rect -1121 883 -1087 917
rect -929 883 -895 917
rect -737 883 -703 917
rect -545 883 -511 917
rect -353 883 -319 917
rect -161 883 -127 917
rect 31 883 65 917
rect 223 883 257 917
rect 415 883 449 917
rect 607 883 641 917
rect 799 883 833 917
rect 991 883 1025 917
rect 1183 883 1217 917
rect 1375 883 1409 917
rect -1409 355 -1375 389
rect -1217 355 -1183 389
rect -1025 355 -991 389
rect -833 355 -799 389
rect -641 355 -607 389
rect -449 355 -415 389
rect -257 355 -223 389
rect -65 355 -31 389
rect 127 355 161 389
rect 319 355 353 389
rect 511 355 545 389
rect 703 355 737 389
rect 895 355 929 389
rect 1087 355 1121 389
rect 1279 355 1313 389
rect -1409 247 -1375 281
rect -1217 247 -1183 281
rect -1025 247 -991 281
rect -833 247 -799 281
rect -641 247 -607 281
rect -449 247 -415 281
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect 511 247 545 281
rect 703 247 737 281
rect 895 247 929 281
rect 1087 247 1121 281
rect 1279 247 1313 281
rect -1313 -281 -1279 -247
rect -1121 -281 -1087 -247
rect -929 -281 -895 -247
rect -737 -281 -703 -247
rect -545 -281 -511 -247
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
rect 415 -281 449 -247
rect 607 -281 641 -247
rect 799 -281 833 -247
rect 991 -281 1025 -247
rect 1183 -281 1217 -247
rect 1375 -281 1409 -247
rect -1313 -389 -1279 -355
rect -1121 -389 -1087 -355
rect -929 -389 -895 -355
rect -737 -389 -703 -355
rect -545 -389 -511 -355
rect -353 -389 -319 -355
rect -161 -389 -127 -355
rect 31 -389 65 -355
rect 223 -389 257 -355
rect 415 -389 449 -355
rect 607 -389 641 -355
rect 799 -389 833 -355
rect 991 -389 1025 -355
rect 1183 -389 1217 -355
rect 1375 -389 1409 -355
rect -1409 -917 -1375 -883
rect -1217 -917 -1183 -883
rect -1025 -917 -991 -883
rect -833 -917 -799 -883
rect -641 -917 -607 -883
rect -449 -917 -415 -883
rect -257 -917 -223 -883
rect -65 -917 -31 -883
rect 127 -917 161 -883
rect 319 -917 353 -883
rect 511 -917 545 -883
rect 703 -917 737 -883
rect 895 -917 929 -883
rect 1087 -917 1121 -883
rect 1279 -917 1313 -883
<< locali >>
rect -1571 985 -1475 1019
rect 1475 985 1571 1019
rect -1571 923 -1537 985
rect 1537 923 1571 985
rect -1329 883 -1313 917
rect -1279 883 -1263 917
rect -1137 883 -1121 917
rect -1087 883 -1071 917
rect -945 883 -929 917
rect -895 883 -879 917
rect -753 883 -737 917
rect -703 883 -687 917
rect -561 883 -545 917
rect -511 883 -495 917
rect -369 883 -353 917
rect -319 883 -303 917
rect -177 883 -161 917
rect -127 883 -111 917
rect 15 883 31 917
rect 65 883 81 917
rect 207 883 223 917
rect 257 883 273 917
rect 399 883 415 917
rect 449 883 465 917
rect 591 883 607 917
rect 641 883 657 917
rect 783 883 799 917
rect 833 883 849 917
rect 975 883 991 917
rect 1025 883 1041 917
rect 1167 883 1183 917
rect 1217 883 1233 917
rect 1359 883 1375 917
rect 1409 883 1425 917
rect -1457 824 -1423 840
rect -1457 432 -1423 448
rect -1361 824 -1327 840
rect -1361 432 -1327 448
rect -1265 824 -1231 840
rect -1265 432 -1231 448
rect -1169 824 -1135 840
rect -1169 432 -1135 448
rect -1073 824 -1039 840
rect -1073 432 -1039 448
rect -977 824 -943 840
rect -977 432 -943 448
rect -881 824 -847 840
rect -881 432 -847 448
rect -785 824 -751 840
rect -785 432 -751 448
rect -689 824 -655 840
rect -689 432 -655 448
rect -593 824 -559 840
rect -593 432 -559 448
rect -497 824 -463 840
rect -497 432 -463 448
rect -401 824 -367 840
rect -401 432 -367 448
rect -305 824 -271 840
rect -305 432 -271 448
rect -209 824 -175 840
rect -209 432 -175 448
rect -113 824 -79 840
rect -113 432 -79 448
rect -17 824 17 840
rect -17 432 17 448
rect 79 824 113 840
rect 79 432 113 448
rect 175 824 209 840
rect 175 432 209 448
rect 271 824 305 840
rect 271 432 305 448
rect 367 824 401 840
rect 367 432 401 448
rect 463 824 497 840
rect 463 432 497 448
rect 559 824 593 840
rect 559 432 593 448
rect 655 824 689 840
rect 655 432 689 448
rect 751 824 785 840
rect 751 432 785 448
rect 847 824 881 840
rect 847 432 881 448
rect 943 824 977 840
rect 943 432 977 448
rect 1039 824 1073 840
rect 1039 432 1073 448
rect 1135 824 1169 840
rect 1135 432 1169 448
rect 1231 824 1265 840
rect 1231 432 1265 448
rect 1327 824 1361 840
rect 1327 432 1361 448
rect 1423 824 1457 840
rect 1423 432 1457 448
rect -1425 355 -1409 389
rect -1375 355 -1359 389
rect -1233 355 -1217 389
rect -1183 355 -1167 389
rect -1041 355 -1025 389
rect -991 355 -975 389
rect -849 355 -833 389
rect -799 355 -783 389
rect -657 355 -641 389
rect -607 355 -591 389
rect -465 355 -449 389
rect -415 355 -399 389
rect -273 355 -257 389
rect -223 355 -207 389
rect -81 355 -65 389
rect -31 355 -15 389
rect 111 355 127 389
rect 161 355 177 389
rect 303 355 319 389
rect 353 355 369 389
rect 495 355 511 389
rect 545 355 561 389
rect 687 355 703 389
rect 737 355 753 389
rect 879 355 895 389
rect 929 355 945 389
rect 1071 355 1087 389
rect 1121 355 1137 389
rect 1263 355 1279 389
rect 1313 355 1329 389
rect -1425 247 -1409 281
rect -1375 247 -1359 281
rect -1233 247 -1217 281
rect -1183 247 -1167 281
rect -1041 247 -1025 281
rect -991 247 -975 281
rect -849 247 -833 281
rect -799 247 -783 281
rect -657 247 -641 281
rect -607 247 -591 281
rect -465 247 -449 281
rect -415 247 -399 281
rect -273 247 -257 281
rect -223 247 -207 281
rect -81 247 -65 281
rect -31 247 -15 281
rect 111 247 127 281
rect 161 247 177 281
rect 303 247 319 281
rect 353 247 369 281
rect 495 247 511 281
rect 545 247 561 281
rect 687 247 703 281
rect 737 247 753 281
rect 879 247 895 281
rect 929 247 945 281
rect 1071 247 1087 281
rect 1121 247 1137 281
rect 1263 247 1279 281
rect 1313 247 1329 281
rect -1457 188 -1423 204
rect -1457 -204 -1423 -188
rect -1361 188 -1327 204
rect -1361 -204 -1327 -188
rect -1265 188 -1231 204
rect -1265 -204 -1231 -188
rect -1169 188 -1135 204
rect -1169 -204 -1135 -188
rect -1073 188 -1039 204
rect -1073 -204 -1039 -188
rect -977 188 -943 204
rect -977 -204 -943 -188
rect -881 188 -847 204
rect -881 -204 -847 -188
rect -785 188 -751 204
rect -785 -204 -751 -188
rect -689 188 -655 204
rect -689 -204 -655 -188
rect -593 188 -559 204
rect -593 -204 -559 -188
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect 559 188 593 204
rect 559 -204 593 -188
rect 655 188 689 204
rect 655 -204 689 -188
rect 751 188 785 204
rect 751 -204 785 -188
rect 847 188 881 204
rect 847 -204 881 -188
rect 943 188 977 204
rect 943 -204 977 -188
rect 1039 188 1073 204
rect 1039 -204 1073 -188
rect 1135 188 1169 204
rect 1135 -204 1169 -188
rect 1231 188 1265 204
rect 1231 -204 1265 -188
rect 1327 188 1361 204
rect 1327 -204 1361 -188
rect 1423 188 1457 204
rect 1423 -204 1457 -188
rect -1329 -281 -1313 -247
rect -1279 -281 -1263 -247
rect -1137 -281 -1121 -247
rect -1087 -281 -1071 -247
rect -945 -281 -929 -247
rect -895 -281 -879 -247
rect -753 -281 -737 -247
rect -703 -281 -687 -247
rect -561 -281 -545 -247
rect -511 -281 -495 -247
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 207 -281 223 -247
rect 257 -281 273 -247
rect 399 -281 415 -247
rect 449 -281 465 -247
rect 591 -281 607 -247
rect 641 -281 657 -247
rect 783 -281 799 -247
rect 833 -281 849 -247
rect 975 -281 991 -247
rect 1025 -281 1041 -247
rect 1167 -281 1183 -247
rect 1217 -281 1233 -247
rect 1359 -281 1375 -247
rect 1409 -281 1425 -247
rect -1329 -389 -1313 -355
rect -1279 -389 -1263 -355
rect -1137 -389 -1121 -355
rect -1087 -389 -1071 -355
rect -945 -389 -929 -355
rect -895 -389 -879 -355
rect -753 -389 -737 -355
rect -703 -389 -687 -355
rect -561 -389 -545 -355
rect -511 -389 -495 -355
rect -369 -389 -353 -355
rect -319 -389 -303 -355
rect -177 -389 -161 -355
rect -127 -389 -111 -355
rect 15 -389 31 -355
rect 65 -389 81 -355
rect 207 -389 223 -355
rect 257 -389 273 -355
rect 399 -389 415 -355
rect 449 -389 465 -355
rect 591 -389 607 -355
rect 641 -389 657 -355
rect 783 -389 799 -355
rect 833 -389 849 -355
rect 975 -389 991 -355
rect 1025 -389 1041 -355
rect 1167 -389 1183 -355
rect 1217 -389 1233 -355
rect 1359 -389 1375 -355
rect 1409 -389 1425 -355
rect -1457 -448 -1423 -432
rect -1457 -840 -1423 -824
rect -1361 -448 -1327 -432
rect -1361 -840 -1327 -824
rect -1265 -448 -1231 -432
rect -1265 -840 -1231 -824
rect -1169 -448 -1135 -432
rect -1169 -840 -1135 -824
rect -1073 -448 -1039 -432
rect -1073 -840 -1039 -824
rect -977 -448 -943 -432
rect -977 -840 -943 -824
rect -881 -448 -847 -432
rect -881 -840 -847 -824
rect -785 -448 -751 -432
rect -785 -840 -751 -824
rect -689 -448 -655 -432
rect -689 -840 -655 -824
rect -593 -448 -559 -432
rect -593 -840 -559 -824
rect -497 -448 -463 -432
rect -497 -840 -463 -824
rect -401 -448 -367 -432
rect -401 -840 -367 -824
rect -305 -448 -271 -432
rect -305 -840 -271 -824
rect -209 -448 -175 -432
rect -209 -840 -175 -824
rect -113 -448 -79 -432
rect -113 -840 -79 -824
rect -17 -448 17 -432
rect -17 -840 17 -824
rect 79 -448 113 -432
rect 79 -840 113 -824
rect 175 -448 209 -432
rect 175 -840 209 -824
rect 271 -448 305 -432
rect 271 -840 305 -824
rect 367 -448 401 -432
rect 367 -840 401 -824
rect 463 -448 497 -432
rect 463 -840 497 -824
rect 559 -448 593 -432
rect 559 -840 593 -824
rect 655 -448 689 -432
rect 655 -840 689 -824
rect 751 -448 785 -432
rect 751 -840 785 -824
rect 847 -448 881 -432
rect 847 -840 881 -824
rect 943 -448 977 -432
rect 943 -840 977 -824
rect 1039 -448 1073 -432
rect 1039 -840 1073 -824
rect 1135 -448 1169 -432
rect 1135 -840 1169 -824
rect 1231 -448 1265 -432
rect 1231 -840 1265 -824
rect 1327 -448 1361 -432
rect 1327 -840 1361 -824
rect 1423 -448 1457 -432
rect 1423 -840 1457 -824
rect -1425 -917 -1409 -883
rect -1375 -917 -1359 -883
rect -1233 -917 -1217 -883
rect -1183 -917 -1167 -883
rect -1041 -917 -1025 -883
rect -991 -917 -975 -883
rect -849 -917 -833 -883
rect -799 -917 -783 -883
rect -657 -917 -641 -883
rect -607 -917 -591 -883
rect -465 -917 -449 -883
rect -415 -917 -399 -883
rect -273 -917 -257 -883
rect -223 -917 -207 -883
rect -81 -917 -65 -883
rect -31 -917 -15 -883
rect 111 -917 127 -883
rect 161 -917 177 -883
rect 303 -917 319 -883
rect 353 -917 369 -883
rect 495 -917 511 -883
rect 545 -917 561 -883
rect 687 -917 703 -883
rect 737 -917 753 -883
rect 879 -917 895 -883
rect 929 -917 945 -883
rect 1071 -917 1087 -883
rect 1121 -917 1137 -883
rect 1263 -917 1279 -883
rect 1313 -917 1329 -883
rect -1571 -985 -1537 -923
rect 1537 -985 1571 -923
rect -1571 -1019 -1475 -985
rect 1475 -1019 1571 -985
<< viali >>
rect -1313 883 -1279 917
rect -1121 883 -1087 917
rect -929 883 -895 917
rect -737 883 -703 917
rect -545 883 -511 917
rect -353 883 -319 917
rect -161 883 -127 917
rect 31 883 65 917
rect 223 883 257 917
rect 415 883 449 917
rect 607 883 641 917
rect 799 883 833 917
rect 991 883 1025 917
rect 1183 883 1217 917
rect 1375 883 1409 917
rect -1457 448 -1423 824
rect -1361 448 -1327 824
rect -1265 448 -1231 824
rect -1169 448 -1135 824
rect -1073 448 -1039 824
rect -977 448 -943 824
rect -881 448 -847 824
rect -785 448 -751 824
rect -689 448 -655 824
rect -593 448 -559 824
rect -497 448 -463 824
rect -401 448 -367 824
rect -305 448 -271 824
rect -209 448 -175 824
rect -113 448 -79 824
rect -17 448 17 824
rect 79 448 113 824
rect 175 448 209 824
rect 271 448 305 824
rect 367 448 401 824
rect 463 448 497 824
rect 559 448 593 824
rect 655 448 689 824
rect 751 448 785 824
rect 847 448 881 824
rect 943 448 977 824
rect 1039 448 1073 824
rect 1135 448 1169 824
rect 1231 448 1265 824
rect 1327 448 1361 824
rect 1423 448 1457 824
rect -1409 355 -1375 389
rect -1217 355 -1183 389
rect -1025 355 -991 389
rect -833 355 -799 389
rect -641 355 -607 389
rect -449 355 -415 389
rect -257 355 -223 389
rect -65 355 -31 389
rect 127 355 161 389
rect 319 355 353 389
rect 511 355 545 389
rect 703 355 737 389
rect 895 355 929 389
rect 1087 355 1121 389
rect 1279 355 1313 389
rect -1409 247 -1375 281
rect -1217 247 -1183 281
rect -1025 247 -991 281
rect -833 247 -799 281
rect -641 247 -607 281
rect -449 247 -415 281
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect 511 247 545 281
rect 703 247 737 281
rect 895 247 929 281
rect 1087 247 1121 281
rect 1279 247 1313 281
rect -1457 -188 -1423 188
rect -1361 -188 -1327 188
rect -1265 -188 -1231 188
rect -1169 -188 -1135 188
rect -1073 -188 -1039 188
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect 1039 -188 1073 188
rect 1135 -188 1169 188
rect 1231 -188 1265 188
rect 1327 -188 1361 188
rect 1423 -188 1457 188
rect -1313 -281 -1279 -247
rect -1121 -281 -1087 -247
rect -929 -281 -895 -247
rect -737 -281 -703 -247
rect -545 -281 -511 -247
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
rect 415 -281 449 -247
rect 607 -281 641 -247
rect 799 -281 833 -247
rect 991 -281 1025 -247
rect 1183 -281 1217 -247
rect 1375 -281 1409 -247
rect -1313 -389 -1279 -355
rect -1121 -389 -1087 -355
rect -929 -389 -895 -355
rect -737 -389 -703 -355
rect -545 -389 -511 -355
rect -353 -389 -319 -355
rect -161 -389 -127 -355
rect 31 -389 65 -355
rect 223 -389 257 -355
rect 415 -389 449 -355
rect 607 -389 641 -355
rect 799 -389 833 -355
rect 991 -389 1025 -355
rect 1183 -389 1217 -355
rect 1375 -389 1409 -355
rect -1457 -824 -1423 -448
rect -1361 -824 -1327 -448
rect -1265 -824 -1231 -448
rect -1169 -824 -1135 -448
rect -1073 -824 -1039 -448
rect -977 -824 -943 -448
rect -881 -824 -847 -448
rect -785 -824 -751 -448
rect -689 -824 -655 -448
rect -593 -824 -559 -448
rect -497 -824 -463 -448
rect -401 -824 -367 -448
rect -305 -824 -271 -448
rect -209 -824 -175 -448
rect -113 -824 -79 -448
rect -17 -824 17 -448
rect 79 -824 113 -448
rect 175 -824 209 -448
rect 271 -824 305 -448
rect 367 -824 401 -448
rect 463 -824 497 -448
rect 559 -824 593 -448
rect 655 -824 689 -448
rect 751 -824 785 -448
rect 847 -824 881 -448
rect 943 -824 977 -448
rect 1039 -824 1073 -448
rect 1135 -824 1169 -448
rect 1231 -824 1265 -448
rect 1327 -824 1361 -448
rect 1423 -824 1457 -448
rect -1409 -917 -1375 -883
rect -1217 -917 -1183 -883
rect -1025 -917 -991 -883
rect -833 -917 -799 -883
rect -641 -917 -607 -883
rect -449 -917 -415 -883
rect -257 -917 -223 -883
rect -65 -917 -31 -883
rect 127 -917 161 -883
rect 319 -917 353 -883
rect 511 -917 545 -883
rect 703 -917 737 -883
rect 895 -917 929 -883
rect 1087 -917 1121 -883
rect 1279 -917 1313 -883
<< metal1 >>
rect -1325 917 -1267 923
rect -1325 883 -1313 917
rect -1279 883 -1267 917
rect -1325 877 -1267 883
rect -1133 917 -1075 923
rect -1133 883 -1121 917
rect -1087 883 -1075 917
rect -1133 877 -1075 883
rect -941 917 -883 923
rect -941 883 -929 917
rect -895 883 -883 917
rect -941 877 -883 883
rect -749 917 -691 923
rect -749 883 -737 917
rect -703 883 -691 917
rect -749 877 -691 883
rect -557 917 -499 923
rect -557 883 -545 917
rect -511 883 -499 917
rect -557 877 -499 883
rect -365 917 -307 923
rect -365 883 -353 917
rect -319 883 -307 917
rect -365 877 -307 883
rect -173 917 -115 923
rect -173 883 -161 917
rect -127 883 -115 917
rect -173 877 -115 883
rect 19 917 77 923
rect 19 883 31 917
rect 65 883 77 917
rect 19 877 77 883
rect 211 917 269 923
rect 211 883 223 917
rect 257 883 269 917
rect 211 877 269 883
rect 403 917 461 923
rect 403 883 415 917
rect 449 883 461 917
rect 403 877 461 883
rect 595 917 653 923
rect 595 883 607 917
rect 641 883 653 917
rect 595 877 653 883
rect 787 917 845 923
rect 787 883 799 917
rect 833 883 845 917
rect 787 877 845 883
rect 979 917 1037 923
rect 979 883 991 917
rect 1025 883 1037 917
rect 979 877 1037 883
rect 1171 917 1229 923
rect 1171 883 1183 917
rect 1217 883 1229 917
rect 1171 877 1229 883
rect 1363 917 1421 923
rect 1363 883 1375 917
rect 1409 883 1421 917
rect 1363 877 1421 883
rect -1463 824 -1417 836
rect -1463 448 -1457 824
rect -1423 448 -1417 824
rect -1463 436 -1417 448
rect -1367 824 -1321 836
rect -1367 448 -1361 824
rect -1327 448 -1321 824
rect -1367 436 -1321 448
rect -1271 824 -1225 836
rect -1271 448 -1265 824
rect -1231 448 -1225 824
rect -1271 436 -1225 448
rect -1175 824 -1129 836
rect -1175 448 -1169 824
rect -1135 448 -1129 824
rect -1175 436 -1129 448
rect -1079 824 -1033 836
rect -1079 448 -1073 824
rect -1039 448 -1033 824
rect -1079 436 -1033 448
rect -983 824 -937 836
rect -983 448 -977 824
rect -943 448 -937 824
rect -983 436 -937 448
rect -887 824 -841 836
rect -887 448 -881 824
rect -847 448 -841 824
rect -887 436 -841 448
rect -791 824 -745 836
rect -791 448 -785 824
rect -751 448 -745 824
rect -791 436 -745 448
rect -695 824 -649 836
rect -695 448 -689 824
rect -655 448 -649 824
rect -695 436 -649 448
rect -599 824 -553 836
rect -599 448 -593 824
rect -559 448 -553 824
rect -599 436 -553 448
rect -503 824 -457 836
rect -503 448 -497 824
rect -463 448 -457 824
rect -503 436 -457 448
rect -407 824 -361 836
rect -407 448 -401 824
rect -367 448 -361 824
rect -407 436 -361 448
rect -311 824 -265 836
rect -311 448 -305 824
rect -271 448 -265 824
rect -311 436 -265 448
rect -215 824 -169 836
rect -215 448 -209 824
rect -175 448 -169 824
rect -215 436 -169 448
rect -119 824 -73 836
rect -119 448 -113 824
rect -79 448 -73 824
rect -119 436 -73 448
rect -23 824 23 836
rect -23 448 -17 824
rect 17 448 23 824
rect -23 436 23 448
rect 73 824 119 836
rect 73 448 79 824
rect 113 448 119 824
rect 73 436 119 448
rect 169 824 215 836
rect 169 448 175 824
rect 209 448 215 824
rect 169 436 215 448
rect 265 824 311 836
rect 265 448 271 824
rect 305 448 311 824
rect 265 436 311 448
rect 361 824 407 836
rect 361 448 367 824
rect 401 448 407 824
rect 361 436 407 448
rect 457 824 503 836
rect 457 448 463 824
rect 497 448 503 824
rect 457 436 503 448
rect 553 824 599 836
rect 553 448 559 824
rect 593 448 599 824
rect 553 436 599 448
rect 649 824 695 836
rect 649 448 655 824
rect 689 448 695 824
rect 649 436 695 448
rect 745 824 791 836
rect 745 448 751 824
rect 785 448 791 824
rect 745 436 791 448
rect 841 824 887 836
rect 841 448 847 824
rect 881 448 887 824
rect 841 436 887 448
rect 937 824 983 836
rect 937 448 943 824
rect 977 448 983 824
rect 937 436 983 448
rect 1033 824 1079 836
rect 1033 448 1039 824
rect 1073 448 1079 824
rect 1033 436 1079 448
rect 1129 824 1175 836
rect 1129 448 1135 824
rect 1169 448 1175 824
rect 1129 436 1175 448
rect 1225 824 1271 836
rect 1225 448 1231 824
rect 1265 448 1271 824
rect 1225 436 1271 448
rect 1321 824 1367 836
rect 1321 448 1327 824
rect 1361 448 1367 824
rect 1321 436 1367 448
rect 1417 824 1463 836
rect 1417 448 1423 824
rect 1457 448 1463 824
rect 1417 436 1463 448
rect -1421 389 -1363 395
rect -1421 355 -1409 389
rect -1375 355 -1363 389
rect -1421 349 -1363 355
rect -1229 389 -1171 395
rect -1229 355 -1217 389
rect -1183 355 -1171 389
rect -1229 349 -1171 355
rect -1037 389 -979 395
rect -1037 355 -1025 389
rect -991 355 -979 389
rect -1037 349 -979 355
rect -845 389 -787 395
rect -845 355 -833 389
rect -799 355 -787 389
rect -845 349 -787 355
rect -653 389 -595 395
rect -653 355 -641 389
rect -607 355 -595 389
rect -653 349 -595 355
rect -461 389 -403 395
rect -461 355 -449 389
rect -415 355 -403 389
rect -461 349 -403 355
rect -269 389 -211 395
rect -269 355 -257 389
rect -223 355 -211 389
rect -269 349 -211 355
rect -77 389 -19 395
rect -77 355 -65 389
rect -31 355 -19 389
rect -77 349 -19 355
rect 115 389 173 395
rect 115 355 127 389
rect 161 355 173 389
rect 115 349 173 355
rect 307 389 365 395
rect 307 355 319 389
rect 353 355 365 389
rect 307 349 365 355
rect 499 389 557 395
rect 499 355 511 389
rect 545 355 557 389
rect 499 349 557 355
rect 691 389 749 395
rect 691 355 703 389
rect 737 355 749 389
rect 691 349 749 355
rect 883 389 941 395
rect 883 355 895 389
rect 929 355 941 389
rect 883 349 941 355
rect 1075 389 1133 395
rect 1075 355 1087 389
rect 1121 355 1133 389
rect 1075 349 1133 355
rect 1267 389 1325 395
rect 1267 355 1279 389
rect 1313 355 1325 389
rect 1267 349 1325 355
rect -1421 281 -1363 287
rect -1421 247 -1409 281
rect -1375 247 -1363 281
rect -1421 241 -1363 247
rect -1229 281 -1171 287
rect -1229 247 -1217 281
rect -1183 247 -1171 281
rect -1229 241 -1171 247
rect -1037 281 -979 287
rect -1037 247 -1025 281
rect -991 247 -979 281
rect -1037 241 -979 247
rect -845 281 -787 287
rect -845 247 -833 281
rect -799 247 -787 281
rect -845 241 -787 247
rect -653 281 -595 287
rect -653 247 -641 281
rect -607 247 -595 281
rect -653 241 -595 247
rect -461 281 -403 287
rect -461 247 -449 281
rect -415 247 -403 281
rect -461 241 -403 247
rect -269 281 -211 287
rect -269 247 -257 281
rect -223 247 -211 281
rect -269 241 -211 247
rect -77 281 -19 287
rect -77 247 -65 281
rect -31 247 -19 281
rect -77 241 -19 247
rect 115 281 173 287
rect 115 247 127 281
rect 161 247 173 281
rect 115 241 173 247
rect 307 281 365 287
rect 307 247 319 281
rect 353 247 365 281
rect 307 241 365 247
rect 499 281 557 287
rect 499 247 511 281
rect 545 247 557 281
rect 499 241 557 247
rect 691 281 749 287
rect 691 247 703 281
rect 737 247 749 281
rect 691 241 749 247
rect 883 281 941 287
rect 883 247 895 281
rect 929 247 941 281
rect 883 241 941 247
rect 1075 281 1133 287
rect 1075 247 1087 281
rect 1121 247 1133 281
rect 1075 241 1133 247
rect 1267 281 1325 287
rect 1267 247 1279 281
rect 1313 247 1325 281
rect 1267 241 1325 247
rect -1463 188 -1417 200
rect -1463 -188 -1457 188
rect -1423 -188 -1417 188
rect -1463 -200 -1417 -188
rect -1367 188 -1321 200
rect -1367 -188 -1361 188
rect -1327 -188 -1321 188
rect -1367 -200 -1321 -188
rect -1271 188 -1225 200
rect -1271 -188 -1265 188
rect -1231 -188 -1225 188
rect -1271 -200 -1225 -188
rect -1175 188 -1129 200
rect -1175 -188 -1169 188
rect -1135 -188 -1129 188
rect -1175 -200 -1129 -188
rect -1079 188 -1033 200
rect -1079 -188 -1073 188
rect -1039 -188 -1033 188
rect -1079 -200 -1033 -188
rect -983 188 -937 200
rect -983 -188 -977 188
rect -943 -188 -937 188
rect -983 -200 -937 -188
rect -887 188 -841 200
rect -887 -188 -881 188
rect -847 -188 -841 188
rect -887 -200 -841 -188
rect -791 188 -745 200
rect -791 -188 -785 188
rect -751 -188 -745 188
rect -791 -200 -745 -188
rect -695 188 -649 200
rect -695 -188 -689 188
rect -655 -188 -649 188
rect -695 -200 -649 -188
rect -599 188 -553 200
rect -599 -188 -593 188
rect -559 -188 -553 188
rect -599 -200 -553 -188
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect 553 188 599 200
rect 553 -188 559 188
rect 593 -188 599 188
rect 553 -200 599 -188
rect 649 188 695 200
rect 649 -188 655 188
rect 689 -188 695 188
rect 649 -200 695 -188
rect 745 188 791 200
rect 745 -188 751 188
rect 785 -188 791 188
rect 745 -200 791 -188
rect 841 188 887 200
rect 841 -188 847 188
rect 881 -188 887 188
rect 841 -200 887 -188
rect 937 188 983 200
rect 937 -188 943 188
rect 977 -188 983 188
rect 937 -200 983 -188
rect 1033 188 1079 200
rect 1033 -188 1039 188
rect 1073 -188 1079 188
rect 1033 -200 1079 -188
rect 1129 188 1175 200
rect 1129 -188 1135 188
rect 1169 -188 1175 188
rect 1129 -200 1175 -188
rect 1225 188 1271 200
rect 1225 -188 1231 188
rect 1265 -188 1271 188
rect 1225 -200 1271 -188
rect 1321 188 1367 200
rect 1321 -188 1327 188
rect 1361 -188 1367 188
rect 1321 -200 1367 -188
rect 1417 188 1463 200
rect 1417 -188 1423 188
rect 1457 -188 1463 188
rect 1417 -200 1463 -188
rect -1325 -247 -1267 -241
rect -1325 -281 -1313 -247
rect -1279 -281 -1267 -247
rect -1325 -287 -1267 -281
rect -1133 -247 -1075 -241
rect -1133 -281 -1121 -247
rect -1087 -281 -1075 -247
rect -1133 -287 -1075 -281
rect -941 -247 -883 -241
rect -941 -281 -929 -247
rect -895 -281 -883 -247
rect -941 -287 -883 -281
rect -749 -247 -691 -241
rect -749 -281 -737 -247
rect -703 -281 -691 -247
rect -749 -287 -691 -281
rect -557 -247 -499 -241
rect -557 -281 -545 -247
rect -511 -281 -499 -247
rect -557 -287 -499 -281
rect -365 -247 -307 -241
rect -365 -281 -353 -247
rect -319 -281 -307 -247
rect -365 -287 -307 -281
rect -173 -247 -115 -241
rect -173 -281 -161 -247
rect -127 -281 -115 -247
rect -173 -287 -115 -281
rect 19 -247 77 -241
rect 19 -281 31 -247
rect 65 -281 77 -247
rect 19 -287 77 -281
rect 211 -247 269 -241
rect 211 -281 223 -247
rect 257 -281 269 -247
rect 211 -287 269 -281
rect 403 -247 461 -241
rect 403 -281 415 -247
rect 449 -281 461 -247
rect 403 -287 461 -281
rect 595 -247 653 -241
rect 595 -281 607 -247
rect 641 -281 653 -247
rect 595 -287 653 -281
rect 787 -247 845 -241
rect 787 -281 799 -247
rect 833 -281 845 -247
rect 787 -287 845 -281
rect 979 -247 1037 -241
rect 979 -281 991 -247
rect 1025 -281 1037 -247
rect 979 -287 1037 -281
rect 1171 -247 1229 -241
rect 1171 -281 1183 -247
rect 1217 -281 1229 -247
rect 1171 -287 1229 -281
rect 1363 -247 1421 -241
rect 1363 -281 1375 -247
rect 1409 -281 1421 -247
rect 1363 -287 1421 -281
rect -1325 -355 -1267 -349
rect -1325 -389 -1313 -355
rect -1279 -389 -1267 -355
rect -1325 -395 -1267 -389
rect -1133 -355 -1075 -349
rect -1133 -389 -1121 -355
rect -1087 -389 -1075 -355
rect -1133 -395 -1075 -389
rect -941 -355 -883 -349
rect -941 -389 -929 -355
rect -895 -389 -883 -355
rect -941 -395 -883 -389
rect -749 -355 -691 -349
rect -749 -389 -737 -355
rect -703 -389 -691 -355
rect -749 -395 -691 -389
rect -557 -355 -499 -349
rect -557 -389 -545 -355
rect -511 -389 -499 -355
rect -557 -395 -499 -389
rect -365 -355 -307 -349
rect -365 -389 -353 -355
rect -319 -389 -307 -355
rect -365 -395 -307 -389
rect -173 -355 -115 -349
rect -173 -389 -161 -355
rect -127 -389 -115 -355
rect -173 -395 -115 -389
rect 19 -355 77 -349
rect 19 -389 31 -355
rect 65 -389 77 -355
rect 19 -395 77 -389
rect 211 -355 269 -349
rect 211 -389 223 -355
rect 257 -389 269 -355
rect 211 -395 269 -389
rect 403 -355 461 -349
rect 403 -389 415 -355
rect 449 -389 461 -355
rect 403 -395 461 -389
rect 595 -355 653 -349
rect 595 -389 607 -355
rect 641 -389 653 -355
rect 595 -395 653 -389
rect 787 -355 845 -349
rect 787 -389 799 -355
rect 833 -389 845 -355
rect 787 -395 845 -389
rect 979 -355 1037 -349
rect 979 -389 991 -355
rect 1025 -389 1037 -355
rect 979 -395 1037 -389
rect 1171 -355 1229 -349
rect 1171 -389 1183 -355
rect 1217 -389 1229 -355
rect 1171 -395 1229 -389
rect 1363 -355 1421 -349
rect 1363 -389 1375 -355
rect 1409 -389 1421 -355
rect 1363 -395 1421 -389
rect -1463 -448 -1417 -436
rect -1463 -824 -1457 -448
rect -1423 -824 -1417 -448
rect -1463 -836 -1417 -824
rect -1367 -448 -1321 -436
rect -1367 -824 -1361 -448
rect -1327 -824 -1321 -448
rect -1367 -836 -1321 -824
rect -1271 -448 -1225 -436
rect -1271 -824 -1265 -448
rect -1231 -824 -1225 -448
rect -1271 -836 -1225 -824
rect -1175 -448 -1129 -436
rect -1175 -824 -1169 -448
rect -1135 -824 -1129 -448
rect -1175 -836 -1129 -824
rect -1079 -448 -1033 -436
rect -1079 -824 -1073 -448
rect -1039 -824 -1033 -448
rect -1079 -836 -1033 -824
rect -983 -448 -937 -436
rect -983 -824 -977 -448
rect -943 -824 -937 -448
rect -983 -836 -937 -824
rect -887 -448 -841 -436
rect -887 -824 -881 -448
rect -847 -824 -841 -448
rect -887 -836 -841 -824
rect -791 -448 -745 -436
rect -791 -824 -785 -448
rect -751 -824 -745 -448
rect -791 -836 -745 -824
rect -695 -448 -649 -436
rect -695 -824 -689 -448
rect -655 -824 -649 -448
rect -695 -836 -649 -824
rect -599 -448 -553 -436
rect -599 -824 -593 -448
rect -559 -824 -553 -448
rect -599 -836 -553 -824
rect -503 -448 -457 -436
rect -503 -824 -497 -448
rect -463 -824 -457 -448
rect -503 -836 -457 -824
rect -407 -448 -361 -436
rect -407 -824 -401 -448
rect -367 -824 -361 -448
rect -407 -836 -361 -824
rect -311 -448 -265 -436
rect -311 -824 -305 -448
rect -271 -824 -265 -448
rect -311 -836 -265 -824
rect -215 -448 -169 -436
rect -215 -824 -209 -448
rect -175 -824 -169 -448
rect -215 -836 -169 -824
rect -119 -448 -73 -436
rect -119 -824 -113 -448
rect -79 -824 -73 -448
rect -119 -836 -73 -824
rect -23 -448 23 -436
rect -23 -824 -17 -448
rect 17 -824 23 -448
rect -23 -836 23 -824
rect 73 -448 119 -436
rect 73 -824 79 -448
rect 113 -824 119 -448
rect 73 -836 119 -824
rect 169 -448 215 -436
rect 169 -824 175 -448
rect 209 -824 215 -448
rect 169 -836 215 -824
rect 265 -448 311 -436
rect 265 -824 271 -448
rect 305 -824 311 -448
rect 265 -836 311 -824
rect 361 -448 407 -436
rect 361 -824 367 -448
rect 401 -824 407 -448
rect 361 -836 407 -824
rect 457 -448 503 -436
rect 457 -824 463 -448
rect 497 -824 503 -448
rect 457 -836 503 -824
rect 553 -448 599 -436
rect 553 -824 559 -448
rect 593 -824 599 -448
rect 553 -836 599 -824
rect 649 -448 695 -436
rect 649 -824 655 -448
rect 689 -824 695 -448
rect 649 -836 695 -824
rect 745 -448 791 -436
rect 745 -824 751 -448
rect 785 -824 791 -448
rect 745 -836 791 -824
rect 841 -448 887 -436
rect 841 -824 847 -448
rect 881 -824 887 -448
rect 841 -836 887 -824
rect 937 -448 983 -436
rect 937 -824 943 -448
rect 977 -824 983 -448
rect 937 -836 983 -824
rect 1033 -448 1079 -436
rect 1033 -824 1039 -448
rect 1073 -824 1079 -448
rect 1033 -836 1079 -824
rect 1129 -448 1175 -436
rect 1129 -824 1135 -448
rect 1169 -824 1175 -448
rect 1129 -836 1175 -824
rect 1225 -448 1271 -436
rect 1225 -824 1231 -448
rect 1265 -824 1271 -448
rect 1225 -836 1271 -824
rect 1321 -448 1367 -436
rect 1321 -824 1327 -448
rect 1361 -824 1367 -448
rect 1321 -836 1367 -824
rect 1417 -448 1463 -436
rect 1417 -824 1423 -448
rect 1457 -824 1463 -448
rect 1417 -836 1463 -824
rect -1421 -883 -1363 -877
rect -1421 -917 -1409 -883
rect -1375 -917 -1363 -883
rect -1421 -923 -1363 -917
rect -1229 -883 -1171 -877
rect -1229 -917 -1217 -883
rect -1183 -917 -1171 -883
rect -1229 -923 -1171 -917
rect -1037 -883 -979 -877
rect -1037 -917 -1025 -883
rect -991 -917 -979 -883
rect -1037 -923 -979 -917
rect -845 -883 -787 -877
rect -845 -917 -833 -883
rect -799 -917 -787 -883
rect -845 -923 -787 -917
rect -653 -883 -595 -877
rect -653 -917 -641 -883
rect -607 -917 -595 -883
rect -653 -923 -595 -917
rect -461 -883 -403 -877
rect -461 -917 -449 -883
rect -415 -917 -403 -883
rect -461 -923 -403 -917
rect -269 -883 -211 -877
rect -269 -917 -257 -883
rect -223 -917 -211 -883
rect -269 -923 -211 -917
rect -77 -883 -19 -877
rect -77 -917 -65 -883
rect -31 -917 -19 -883
rect -77 -923 -19 -917
rect 115 -883 173 -877
rect 115 -917 127 -883
rect 161 -917 173 -883
rect 115 -923 173 -917
rect 307 -883 365 -877
rect 307 -917 319 -883
rect 353 -917 365 -883
rect 307 -923 365 -917
rect 499 -883 557 -877
rect 499 -917 511 -883
rect 545 -917 557 -883
rect 499 -923 557 -917
rect 691 -883 749 -877
rect 691 -917 703 -883
rect 737 -917 749 -883
rect 691 -923 749 -917
rect 883 -883 941 -877
rect 883 -917 895 -883
rect 929 -917 941 -883
rect 883 -923 941 -917
rect 1075 -883 1133 -877
rect 1075 -917 1087 -883
rect 1121 -917 1133 -883
rect 1075 -923 1133 -917
rect 1267 -883 1325 -877
rect 1267 -917 1279 -883
rect 1313 -917 1325 -883
rect 1267 -923 1325 -917
<< properties >>
string FIXED_BBOX -1554 -1002 1554 1002
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 3 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
