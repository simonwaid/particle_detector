magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< nwell >>
rect -10 1380 1100 1390
rect 940 550 1100 1380
rect 172 376 910 442
rect 286 370 316 376
rect 478 370 508 376
rect 670 370 700 376
rect 862 370 892 376
rect 190 -86 220 -80
rect 382 -86 412 -80
rect 574 -86 604 -80
rect 766 -86 796 -80
rect 172 -152 910 -86
rect 172 -260 910 -194
rect 190 -266 220 -260
rect 382 -266 412 -260
rect 574 -266 604 -260
rect 766 -266 796 -260
rect 286 -722 316 -716
rect 478 -722 508 -716
rect 670 -722 700 -716
rect 862 -722 892 -716
rect 172 -788 910 -722
rect 1080 -910 1100 550
<< poly >>
rect 172 426 910 442
rect 172 392 284 426
rect 318 392 476 426
rect 510 392 668 426
rect 702 392 860 426
rect 894 392 910 426
rect 172 376 910 392
rect 286 370 316 376
rect 478 370 508 376
rect 670 370 700 376
rect 862 370 892 376
rect 190 -86 220 -80
rect 382 -86 412 -80
rect 574 -86 604 -80
rect 766 -86 796 -80
rect 172 -102 910 -86
rect 172 -136 188 -102
rect 222 -136 380 -102
rect 414 -136 572 -102
rect 606 -136 764 -102
rect 798 -136 910 -102
rect 172 -152 910 -136
rect 172 -210 910 -194
rect 172 -244 188 -210
rect 222 -244 380 -210
rect 414 -244 572 -210
rect 606 -244 764 -210
rect 798 -244 910 -210
rect 172 -260 910 -244
rect 190 -266 220 -260
rect 382 -266 412 -260
rect 574 -266 604 -260
rect 766 -266 796 -260
rect 286 -722 316 -716
rect 478 -722 508 -716
rect 670 -722 700 -716
rect 862 -722 892 -716
rect 172 -738 910 -722
rect 172 -772 284 -738
rect 318 -772 476 -738
rect 510 -772 668 -738
rect 702 -772 860 -738
rect 894 -772 910 -738
rect 172 -788 910 -772
<< polycont >>
rect 284 392 318 426
rect 476 392 510 426
rect 668 392 702 426
rect 860 392 894 426
rect 188 -136 222 -102
rect 380 -136 414 -102
rect 572 -136 606 -102
rect 764 -136 798 -102
rect 188 -244 222 -210
rect 380 -244 414 -210
rect 572 -244 606 -210
rect 764 -244 798 -210
rect 284 -772 318 -738
rect 476 -772 510 -738
rect 668 -772 702 -738
rect 860 -772 894 -738
<< locali >>
rect 20 520 920 610
rect 172 392 284 426
rect 318 392 476 426
rect 510 392 668 426
rect 702 392 860 426
rect 894 392 910 426
rect 172 -136 188 -102
rect 222 -136 380 -102
rect 414 -136 572 -102
rect 606 -136 764 -102
rect 798 -136 910 -102
rect 172 -244 188 -210
rect 222 -244 380 -210
rect 414 -244 572 -210
rect 606 -244 764 -210
rect 798 -244 910 -210
rect 172 -772 284 -738
rect 318 -772 476 -738
rect 510 -772 668 -738
rect 702 -772 860 -738
rect 894 -772 910 -738
<< viali >>
rect 380 1300 560 1360
rect 284 392 318 426
rect 476 392 510 426
rect 668 392 702 426
rect 860 392 894 426
rect 188 -136 222 -102
rect 380 -136 414 -102
rect 572 -136 606 -102
rect 764 -136 798 -102
rect 188 -244 222 -210
rect 380 -244 414 -210
rect 572 -244 606 -210
rect 764 -244 798 -210
rect 284 -772 318 -738
rect 476 -772 510 -738
rect 668 -772 702 -738
rect 860 -772 894 -738
<< metal1 >>
rect 368 1360 572 1366
rect 368 1300 380 1360
rect 560 1300 572 1360
rect 368 1294 572 1300
rect 40 1210 760 1260
rect 40 730 90 1210
rect 278 994 288 1170
rect 342 994 352 1170
rect 594 994 604 1170
rect 658 994 668 1170
rect 120 768 130 944
rect 184 768 194 944
rect 436 768 446 944
rect 500 768 510 944
rect 752 768 762 944
rect 816 768 826 944
rect 40 680 760 730
rect 40 440 90 680
rect 40 426 910 440
rect 40 392 284 426
rect 318 392 476 426
rect 510 392 668 426
rect 702 392 860 426
rect 894 392 910 426
rect 40 380 910 392
rect 40 -90 90 380
rect 216 170 226 346
rect 280 170 290 346
rect 408 170 418 346
rect 472 170 482 346
rect 600 170 610 346
rect 664 170 674 346
rect 792 170 802 346
rect 856 170 866 346
rect 120 -56 130 120
rect 184 -56 194 120
rect 312 -56 322 120
rect 376 -56 386 120
rect 504 -56 514 120
rect 568 -56 578 120
rect 696 -56 706 120
rect 760 -56 770 120
rect 888 -56 898 120
rect 952 -56 962 120
rect 40 -102 910 -90
rect 40 -136 188 -102
rect 222 -136 380 -102
rect 414 -136 572 -102
rect 606 -136 764 -102
rect 798 -136 910 -102
rect 40 -150 910 -136
rect 40 -200 90 -150
rect 40 -210 910 -200
rect 40 -244 188 -210
rect 222 -244 380 -210
rect 414 -244 572 -210
rect 606 -244 764 -210
rect 798 -244 910 -210
rect 40 -260 910 -244
rect 40 -730 90 -260
rect 216 -466 226 -290
rect 280 -466 290 -290
rect 408 -466 418 -290
rect 472 -466 482 -290
rect 600 -466 610 -290
rect 664 -466 674 -290
rect 792 -466 802 -290
rect 856 -466 866 -290
rect 120 -692 130 -516
rect 184 -692 194 -516
rect 312 -692 322 -516
rect 376 -692 386 -516
rect 504 -692 514 -516
rect 568 -692 578 -516
rect 696 -692 706 -516
rect 760 -692 770 -516
rect 888 -692 898 -516
rect 952 -692 962 -516
rect 40 -738 910 -730
rect 40 -772 284 -738
rect 318 -772 476 -738
rect 510 -772 668 -738
rect 702 -772 860 -738
rect 894 -772 910 -738
rect 40 -790 910 -772
<< via1 >>
rect 380 1300 560 1360
rect 288 994 342 1170
rect 604 994 658 1170
rect 130 768 184 944
rect 446 768 500 944
rect 762 768 816 944
rect 226 170 280 346
rect 418 170 472 346
rect 610 170 664 346
rect 802 170 856 346
rect 130 -56 184 120
rect 322 -56 376 120
rect 514 -56 568 120
rect 706 -56 760 120
rect 898 -56 952 120
rect 226 -466 280 -290
rect 418 -466 472 -290
rect 610 -466 664 -290
rect 802 -466 856 -290
rect 130 -692 184 -516
rect 322 -692 376 -516
rect 514 -692 568 -516
rect 706 -692 760 -516
rect 898 -692 952 -516
<< metal2 >>
rect 380 1360 560 1370
rect 270 1300 380 1350
rect 560 1300 680 1350
rect 270 1170 680 1300
rect 270 1030 288 1170
rect 342 1030 604 1170
rect 288 984 342 994
rect 658 1030 680 1170
rect 604 984 658 994
rect 130 944 184 954
rect 120 768 130 900
rect 446 944 500 954
rect 184 768 446 900
rect 762 944 816 954
rect 500 768 762 900
rect 816 768 1030 900
rect 120 750 1030 768
rect 210 350 870 360
rect 210 346 620 350
rect 210 210 226 346
rect 280 210 418 346
rect 226 160 280 170
rect 472 210 610 346
rect 860 220 870 350
rect 418 160 472 170
rect 664 210 802 220
rect 610 160 664 170
rect 856 210 870 220
rect 802 160 856 170
rect 910 130 1030 750
rect 130 120 184 130
rect 120 -56 130 80
rect 322 120 376 130
rect 184 -56 322 80
rect 514 120 568 130
rect 376 -56 514 80
rect 706 120 760 130
rect 568 -56 706 80
rect 898 120 1030 130
rect 760 -56 898 80
rect 952 -56 1030 120
rect 120 -70 1030 -56
rect 210 -280 870 -270
rect 210 -290 620 -280
rect 210 -420 226 -290
rect 280 -420 418 -290
rect 226 -476 280 -466
rect 472 -420 610 -290
rect 860 -410 870 -280
rect 418 -476 472 -466
rect 664 -420 802 -410
rect 610 -476 664 -466
rect 856 -420 870 -410
rect 802 -476 856 -466
rect 910 -506 1030 -70
rect 130 -516 184 -506
rect 120 -692 130 -560
rect 322 -516 376 -506
rect 184 -692 322 -560
rect 514 -516 568 -506
rect 376 -692 514 -560
rect 706 -516 760 -506
rect 568 -692 706 -560
rect 898 -516 1030 -506
rect 760 -692 898 -560
rect 952 -692 1030 -516
rect 120 -710 1030 -692
<< via2 >>
rect 620 346 860 350
rect 620 220 664 346
rect 664 220 802 346
rect 802 220 856 346
rect 856 220 860 346
rect 620 -290 860 -280
rect 620 -410 664 -290
rect 664 -410 802 -290
rect 802 -410 856 -290
rect 856 -410 860 -290
<< metal3 >>
rect 610 350 870 355
rect 610 220 620 350
rect 860 220 870 350
rect 610 215 870 220
rect 620 -275 860 215
rect 610 -280 870 -275
rect 610 -410 620 -280
rect 860 -410 870 -280
rect 610 -415 870 -410
use sky130_fd_pr__pfet_01v8_PDCJZ5  sky130_fd_pr__pfet_01v8_PDCJZ5_0
timestamp 1654768133
transform 1 0 473 0 1 969
box -483 -419 483 419
use sky130_fd_pr__pfet_01v8_U4PLGH  sky130_fd_pr__pfet_01v8_U4PLGH_0
timestamp 1654768133
transform 1 0 541 0 1 -173
box -551 -737 551 737
<< end >>
