magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< pwell >>
rect 132 2010 870 2076
rect 132 1500 870 1566
rect 132 1392 870 1458
rect 132 882 870 948
<< poly >>
rect 132 2060 870 2076
rect 132 2026 244 2060
rect 278 2026 436 2060
rect 470 2026 628 2060
rect 662 2026 820 2060
rect 854 2026 870 2060
rect 132 2010 870 2026
rect 132 1550 870 1566
rect 132 1516 148 1550
rect 182 1516 340 1550
rect 374 1516 532 1550
rect 566 1516 724 1550
rect 758 1516 870 1550
rect 132 1500 870 1516
rect 132 1442 870 1458
rect 132 1408 148 1442
rect 182 1408 340 1442
rect 374 1408 532 1442
rect 566 1408 724 1442
rect 758 1408 870 1442
rect 132 1392 870 1408
rect 132 932 870 948
rect 132 898 244 932
rect 278 898 436 932
rect 470 898 628 932
rect 662 898 820 932
rect 854 898 870 932
rect 132 882 870 898
<< polycont >>
rect 244 2026 278 2060
rect 436 2026 470 2060
rect 628 2026 662 2060
rect 820 2026 854 2060
rect 148 1516 182 1550
rect 340 1516 374 1550
rect 532 1516 566 1550
rect 724 1516 758 1550
rect 148 1408 182 1442
rect 340 1408 374 1442
rect 532 1408 566 1442
rect 724 1408 758 1442
rect 244 898 278 932
rect 436 898 470 932
rect 628 898 662 932
rect 820 898 854 932
<< locali >>
rect 132 2026 244 2060
rect 278 2026 436 2060
rect 470 2026 628 2060
rect 662 2026 820 2060
rect 854 2026 870 2060
rect 132 1516 148 1550
rect 182 1516 340 1550
rect 374 1516 532 1550
rect 566 1516 724 1550
rect 758 1516 870 1550
rect 132 1408 148 1442
rect 182 1408 340 1442
rect 374 1408 532 1442
rect 566 1408 724 1442
rect 758 1408 870 1442
rect 132 898 244 932
rect 278 898 436 932
rect 470 898 628 932
rect 662 898 820 932
rect 854 898 870 932
<< viali >>
rect 244 2026 278 2060
rect 436 2026 470 2060
rect 628 2026 662 2060
rect 820 2026 854 2060
rect 148 1516 182 1550
rect 340 1516 374 1550
rect 532 1516 566 1550
rect 724 1516 758 1550
rect 148 1408 182 1442
rect 340 1408 374 1442
rect 532 1408 566 1442
rect 724 1408 758 1442
rect 244 898 278 932
rect 436 898 470 932
rect 628 898 662 932
rect 820 898 854 932
rect 330 -30 550 40
<< metal1 >>
rect 0 2060 870 2070
rect 0 2026 244 2060
rect 278 2026 436 2060
rect 470 2026 628 2060
rect 662 2026 820 2060
rect 854 2026 870 2060
rect 0 2020 870 2026
rect 0 1560 50 2020
rect 176 1812 186 1988
rect 240 1812 250 1988
rect 368 1812 378 1988
rect 432 1812 442 1988
rect 560 1812 570 1988
rect 624 1812 634 1988
rect 752 1812 762 1988
rect 816 1812 826 1988
rect 80 1588 90 1764
rect 144 1588 154 1764
rect 272 1588 282 1764
rect 336 1588 346 1764
rect 464 1588 474 1764
rect 528 1588 538 1764
rect 656 1588 666 1764
rect 720 1588 730 1764
rect 848 1588 858 1764
rect 912 1588 922 1764
rect 0 1550 870 1560
rect 0 1516 148 1550
rect 182 1516 340 1550
rect 374 1516 532 1550
rect 566 1516 724 1550
rect 758 1516 870 1550
rect 0 1510 870 1516
rect 0 1450 50 1510
rect 0 1442 870 1450
rect 0 1408 148 1442
rect 182 1408 340 1442
rect 374 1408 532 1442
rect 566 1408 724 1442
rect 758 1408 870 1442
rect 0 1400 870 1408
rect 0 940 50 1400
rect 176 1194 186 1370
rect 240 1194 250 1370
rect 368 1194 378 1370
rect 432 1194 442 1370
rect 560 1194 570 1370
rect 624 1194 634 1370
rect 752 1194 762 1370
rect 816 1194 826 1370
rect 80 970 90 1146
rect 144 970 154 1146
rect 272 970 282 1146
rect 336 970 346 1146
rect 464 970 474 1146
rect 528 970 538 1146
rect 656 970 666 1146
rect 720 970 730 1146
rect 848 970 858 1146
rect 912 970 922 1146
rect 0 932 870 940
rect 0 898 244 932
rect 278 898 436 932
rect 470 898 628 932
rect 662 898 820 932
rect 854 898 870 932
rect 0 890 870 898
rect 0 640 50 890
rect 0 590 720 640
rect 0 130 50 590
rect 238 384 248 560
rect 302 384 312 560
rect 554 384 564 560
rect 618 384 628 560
rect 80 160 90 336
rect 144 160 154 336
rect 396 160 406 336
rect 460 160 470 336
rect 712 160 722 336
rect 776 160 786 336
rect 0 80 720 130
rect 318 40 562 46
rect 318 -30 330 40
rect 550 -30 562 40
rect 318 -36 562 -30
<< via1 >>
rect 186 1812 240 1988
rect 378 1812 432 1988
rect 570 1812 624 1988
rect 762 1812 816 1988
rect 90 1588 144 1764
rect 282 1588 336 1764
rect 474 1588 528 1764
rect 666 1588 720 1764
rect 858 1588 912 1764
rect 186 1194 240 1370
rect 378 1194 432 1370
rect 570 1194 624 1370
rect 762 1194 816 1370
rect 90 970 144 1146
rect 282 970 336 1146
rect 474 970 528 1146
rect 666 970 720 1146
rect 858 970 912 1146
rect 248 384 302 560
rect 564 384 618 560
rect 90 160 144 336
rect 406 160 460 336
rect 722 160 776 336
rect 330 -30 550 40
<< metal2 >>
rect 170 1990 820 2000
rect 170 1988 580 1990
rect 810 1988 820 1990
rect 170 1850 186 1988
rect 240 1850 378 1988
rect 186 1802 240 1812
rect 432 1850 570 1988
rect 378 1802 432 1812
rect 624 1850 762 1860
rect 570 1802 624 1812
rect 816 1850 820 1988
rect 762 1802 816 1812
rect 90 1764 144 1774
rect 80 1588 90 1720
rect 282 1764 336 1774
rect 144 1588 282 1720
rect 474 1764 528 1774
rect 336 1588 474 1720
rect 666 1764 720 1774
rect 528 1588 666 1720
rect 858 1764 912 1774
rect 720 1588 858 1720
rect 912 1588 1030 1720
rect 80 1570 1030 1588
rect 180 1380 820 1390
rect 180 1370 580 1380
rect 810 1370 820 1380
rect 180 1240 186 1370
rect 240 1240 378 1370
rect 186 1184 240 1194
rect 432 1240 570 1370
rect 378 1184 432 1194
rect 624 1240 762 1250
rect 570 1184 624 1194
rect 816 1240 820 1370
rect 762 1184 816 1194
rect 860 1156 1030 1570
rect 90 1146 144 1156
rect 80 970 90 1110
rect 282 1146 336 1156
rect 144 970 282 1110
rect 474 1146 528 1156
rect 336 970 474 1110
rect 666 1146 720 1156
rect 528 970 666 1110
rect 858 1146 1030 1156
rect 720 970 858 1110
rect 912 970 1030 1146
rect 80 960 1030 970
rect 860 580 1030 960
rect 230 560 1030 580
rect 230 430 248 560
rect 302 430 564 560
rect 248 374 302 384
rect 618 430 1030 560
rect 564 374 618 384
rect 90 336 144 346
rect 80 160 90 290
rect 406 336 460 346
rect 144 160 406 290
rect 722 336 776 346
rect 460 160 722 290
rect 776 160 780 290
rect 80 140 780 160
rect 330 40 550 140
rect 330 -40 550 -30
<< via2 >>
rect 580 1988 810 1990
rect 580 1860 624 1988
rect 624 1860 762 1988
rect 762 1860 810 1988
rect 580 1370 810 1380
rect 580 1250 624 1370
rect 624 1250 762 1370
rect 762 1250 810 1370
<< metal3 >>
rect 560 1990 820 2000
rect 560 1860 580 1990
rect 810 1860 820 1990
rect 560 1380 820 1860
rect 560 1250 580 1380
rect 810 1250 820 1380
rect 560 1240 820 1250
use sky130_fd_pr__nfet_01v8_6YE2KS  sky130_fd_pr__nfet_01v8_6YE2KS_0
timestamp 1654760956
transform 1 0 433 0 1 360
box -483 -410 483 410
use sky130_fd_pr__nfet_01v8_QQ8PGA  sky130_fd_pr__nfet_01v8_QQ8PGA_0
timestamp 1654760956
transform 1 0 501 0 1 1479
box -551 -719 551 719
<< end >>
