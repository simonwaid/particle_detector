magic
tech sky130B
magscale 1 2
timestamp 1654097953
<< pwell >>
rect 352 542 514 608
rect 352 32 514 98
<< poly >>
rect 352 592 514 608
rect 352 558 368 592
rect 402 558 514 592
rect 352 542 514 558
rect 352 82 514 98
rect 352 48 464 82
rect 498 48 514 82
rect 352 32 514 48
<< polycont >>
rect 368 558 402 592
rect 464 48 498 82
<< locali >>
rect 352 558 368 592
rect 402 558 514 592
rect 352 48 464 82
rect 498 48 514 82
rect 0 -130 890 -30
<< viali >>
rect 368 558 402 592
rect 464 48 498 82
rect 340 -1510 550 -1440
<< metal1 >>
rect 210 592 660 600
rect 210 558 368 592
rect 402 558 660 592
rect 210 550 660 558
rect 210 90 260 550
rect 396 344 406 520
rect 460 344 470 520
rect 300 120 310 296
rect 364 120 374 296
rect 492 120 502 296
rect 556 120 566 296
rect 610 90 660 550
rect 210 82 660 90
rect 210 48 464 82
rect 498 48 660 82
rect 210 40 660 48
rect 210 -210 260 40
rect 610 -210 660 40
rect 0 -260 890 -210
rect 0 -720 50 -260
rect 248 -468 258 -292
rect 312 -468 322 -292
rect 564 -468 574 -292
rect 628 -468 638 -292
rect 90 -692 100 -516
rect 154 -692 164 -516
rect 406 -692 416 -516
rect 470 -692 480 -516
rect 722 -692 732 -516
rect 786 -692 796 -516
rect 840 -720 890 -260
rect 0 -770 890 -720
rect 0 -830 50 -770
rect 840 -830 890 -770
rect 0 -880 890 -830
rect 0 -1340 50 -880
rect 248 -1086 258 -910
rect 312 -1086 322 -910
rect 564 -1086 574 -910
rect 628 -1086 638 -910
rect 90 -1310 100 -1134
rect 154 -1310 164 -1134
rect 406 -1310 416 -1134
rect 470 -1310 480 -1134
rect 722 -1310 732 -1134
rect 786 -1310 796 -1134
rect 840 -1340 890 -880
rect 0 -1390 890 -1340
rect 328 -1440 562 -1434
rect 328 -1510 340 -1440
rect 550 -1510 562 -1440
rect 328 -1516 562 -1510
<< via1 >>
rect 406 344 460 520
rect 310 120 364 296
rect 502 120 556 296
rect 258 -468 312 -292
rect 574 -468 628 -292
rect 100 -692 154 -516
rect 416 -692 470 -516
rect 732 -692 786 -516
rect 258 -1086 312 -910
rect 574 -1086 628 -910
rect 100 -1310 154 -1134
rect 416 -1310 470 -1134
rect 732 -1310 786 -1134
rect 340 -1510 550 -1440
<< metal2 >>
rect 406 520 460 530
rect 406 334 460 344
rect 310 300 364 306
rect 502 300 556 306
rect 260 296 630 300
rect 260 290 310 296
rect 364 290 502 296
rect 556 290 630 296
rect 260 110 630 120
rect 250 -290 640 -280
rect 250 -292 260 -290
rect 250 -468 258 -292
rect 630 -460 640 -290
rect 312 -468 574 -460
rect 628 -468 640 -460
rect 250 -470 640 -468
rect 258 -478 312 -470
rect 574 -478 628 -470
rect 100 -510 154 -506
rect 416 -510 470 -506
rect 732 -510 786 -506
rect -10 -516 890 -510
rect -10 -692 100 -516
rect 154 -692 416 -516
rect 470 -692 732 -516
rect 786 -692 890 -516
rect -10 -710 890 -692
rect -10 -1130 200 -710
rect 250 -910 640 -900
rect 250 -1086 258 -910
rect 630 -1080 640 -910
rect 312 -1086 574 -1080
rect 628 -1086 640 -1080
rect 250 -1090 640 -1086
rect 258 -1096 312 -1090
rect 574 -1096 628 -1090
rect 416 -1130 470 -1124
rect 680 -1130 890 -710
rect -10 -1134 890 -1130
rect -10 -1310 100 -1134
rect 154 -1310 416 -1134
rect 470 -1310 732 -1134
rect 786 -1310 890 -1134
rect -10 -1320 890 -1310
rect 340 -1440 550 -1320
rect 340 -1520 550 -1510
<< via2 >>
rect 260 120 310 290
rect 310 120 364 290
rect 364 120 502 290
rect 502 120 556 290
rect 556 120 630 290
rect 260 -292 630 -290
rect 260 -460 312 -292
rect 312 -460 574 -292
rect 574 -460 628 -292
rect 628 -460 630 -292
rect 260 -1080 312 -910
rect 312 -1080 574 -910
rect 574 -1080 628 -910
rect 628 -1080 630 -910
<< metal3 >>
rect 250 290 640 295
rect 250 120 260 290
rect 630 120 640 290
rect 250 115 640 120
rect 260 -285 630 115
rect 250 -290 640 -285
rect 250 -460 260 -290
rect 630 -460 640 -290
rect 250 -465 640 -460
rect 260 -905 630 -465
rect 250 -910 640 -905
rect 250 -1080 260 -910
rect 630 -1080 640 -910
rect 250 -1085 640 -1080
use sky130_fd_pr__nfet_01v8_LH2JGW  sky130_fd_pr__nfet_01v8_LH2JGW_0
timestamp 1654097953
transform 1 0 433 0 1 320
box -263 -410 263 410
use sky130_fd_pr__nfet_01v8_MJG2KS  sky130_fd_pr__nfet_01v8_MJG2KS_0
timestamp 1654074216
transform 1 0 443 0 1 -801
box -483 -719 483 719
<< end >>
