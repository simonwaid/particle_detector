magic
tech sky130A
magscale 1 2
timestamp 1645531774
<< nwell >>
rect -6773 127 -6107 1309
rect -5853 127 -5187 1309
rect -4933 127 -4267 1309
rect -4013 127 -3347 1309
rect -3093 127 -2427 1309
rect -2173 127 -1507 1309
rect -1253 127 -587 1309
rect -333 127 333 1309
rect 587 127 1253 1309
rect 1507 127 2173 1309
rect 2427 127 3093 1309
rect 3347 127 4013 1309
rect 4267 127 4933 1309
rect 5187 127 5853 1309
rect 6107 127 6773 1309
rect -6773 -1309 -6107 -127
rect -5853 -1309 -5187 -127
rect -4933 -1309 -4267 -127
rect -4013 -1309 -3347 -127
rect -3093 -1309 -2427 -127
rect -2173 -1309 -1507 -127
rect -1253 -1309 -587 -127
rect -333 -1309 333 -127
rect 587 -1309 1253 -127
rect 1507 -1309 2173 -127
rect 2427 -1309 3093 -127
rect 3347 -1309 4013 -127
rect 4267 -1309 4933 -127
rect 5187 -1309 5853 -127
rect 6107 -1309 6773 -127
<< pwell >>
rect -6883 1309 6883 1419
rect -6883 127 -6773 1309
rect -6107 127 -5853 1309
rect -5187 127 -4933 1309
rect -4267 127 -4013 1309
rect -3347 127 -3093 1309
rect -2427 127 -2173 1309
rect -1507 127 -1253 1309
rect -587 127 -333 1309
rect 333 127 587 1309
rect 1253 127 1507 1309
rect 2173 127 2427 1309
rect 3093 127 3347 1309
rect 4013 127 4267 1309
rect 4933 127 5187 1309
rect 5853 127 6107 1309
rect 6773 127 6883 1309
rect -6883 -127 6883 127
rect -6883 -1309 -6773 -127
rect -6107 -1309 -5853 -127
rect -5187 -1309 -4933 -127
rect -4267 -1309 -4013 -127
rect -3347 -1309 -3093 -127
rect -2427 -1309 -2173 -127
rect -1507 -1309 -1253 -127
rect -587 -1309 -333 -127
rect 333 -1309 587 -127
rect 1253 -1309 1507 -127
rect 2173 -1309 2427 -127
rect 3093 -1309 3347 -127
rect 4013 -1309 4267 -127
rect 4933 -1309 5187 -127
rect 5853 -1309 6107 -127
rect 6773 -1309 6883 -127
rect -6883 -1419 6883 -1309
<< varactor >>
rect -6640 218 -6240 1218
rect -5720 218 -5320 1218
rect -4800 218 -4400 1218
rect -3880 218 -3480 1218
rect -2960 218 -2560 1218
rect -2040 218 -1640 1218
rect -1120 218 -720 1218
rect -200 218 200 1218
rect 720 218 1120 1218
rect 1640 218 2040 1218
rect 2560 218 2960 1218
rect 3480 218 3880 1218
rect 4400 218 4800 1218
rect 5320 218 5720 1218
rect 6240 218 6640 1218
rect -6640 -1218 -6240 -218
rect -5720 -1218 -5320 -218
rect -4800 -1218 -4400 -218
rect -3880 -1218 -3480 -218
rect -2960 -1218 -2560 -218
rect -2040 -1218 -1640 -218
rect -1120 -1218 -720 -218
rect -200 -1218 200 -218
rect 720 -1218 1120 -218
rect 1640 -1218 2040 -218
rect 2560 -1218 2960 -218
rect 3480 -1218 3880 -218
rect 4400 -1218 4800 -218
rect 5320 -1218 5720 -218
rect 6240 -1218 6640 -218
<< psubdiff >>
rect -6847 1349 -6751 1383
rect 6751 1349 6847 1383
rect -6847 1287 -6813 1349
rect 6813 1287 6847 1349
rect -6847 -1349 -6813 -1287
rect 6813 -1349 6847 -1287
rect -6847 -1383 -6751 -1349
rect 6751 -1383 6847 -1349
<< nsubdiff >>
rect -6737 1194 -6640 1218
rect -6737 242 -6725 1194
rect -6691 242 -6640 1194
rect -6737 218 -6640 242
rect -6240 1194 -6143 1218
rect -6240 242 -6189 1194
rect -6155 242 -6143 1194
rect -6240 218 -6143 242
rect -5817 1194 -5720 1218
rect -5817 242 -5805 1194
rect -5771 242 -5720 1194
rect -5817 218 -5720 242
rect -5320 1194 -5223 1218
rect -5320 242 -5269 1194
rect -5235 242 -5223 1194
rect -5320 218 -5223 242
rect -4897 1194 -4800 1218
rect -4897 242 -4885 1194
rect -4851 242 -4800 1194
rect -4897 218 -4800 242
rect -4400 1194 -4303 1218
rect -4400 242 -4349 1194
rect -4315 242 -4303 1194
rect -4400 218 -4303 242
rect -3977 1194 -3880 1218
rect -3977 242 -3965 1194
rect -3931 242 -3880 1194
rect -3977 218 -3880 242
rect -3480 1194 -3383 1218
rect -3480 242 -3429 1194
rect -3395 242 -3383 1194
rect -3480 218 -3383 242
rect -3057 1194 -2960 1218
rect -3057 242 -3045 1194
rect -3011 242 -2960 1194
rect -3057 218 -2960 242
rect -2560 1194 -2463 1218
rect -2560 242 -2509 1194
rect -2475 242 -2463 1194
rect -2560 218 -2463 242
rect -2137 1194 -2040 1218
rect -2137 242 -2125 1194
rect -2091 242 -2040 1194
rect -2137 218 -2040 242
rect -1640 1194 -1543 1218
rect -1640 242 -1589 1194
rect -1555 242 -1543 1194
rect -1640 218 -1543 242
rect -1217 1194 -1120 1218
rect -1217 242 -1205 1194
rect -1171 242 -1120 1194
rect -1217 218 -1120 242
rect -720 1194 -623 1218
rect -720 242 -669 1194
rect -635 242 -623 1194
rect -720 218 -623 242
rect -297 1194 -200 1218
rect -297 242 -285 1194
rect -251 242 -200 1194
rect -297 218 -200 242
rect 200 1194 297 1218
rect 200 242 251 1194
rect 285 242 297 1194
rect 200 218 297 242
rect 623 1194 720 1218
rect 623 242 635 1194
rect 669 242 720 1194
rect 623 218 720 242
rect 1120 1194 1217 1218
rect 1120 242 1171 1194
rect 1205 242 1217 1194
rect 1120 218 1217 242
rect 1543 1194 1640 1218
rect 1543 242 1555 1194
rect 1589 242 1640 1194
rect 1543 218 1640 242
rect 2040 1194 2137 1218
rect 2040 242 2091 1194
rect 2125 242 2137 1194
rect 2040 218 2137 242
rect 2463 1194 2560 1218
rect 2463 242 2475 1194
rect 2509 242 2560 1194
rect 2463 218 2560 242
rect 2960 1194 3057 1218
rect 2960 242 3011 1194
rect 3045 242 3057 1194
rect 2960 218 3057 242
rect 3383 1194 3480 1218
rect 3383 242 3395 1194
rect 3429 242 3480 1194
rect 3383 218 3480 242
rect 3880 1194 3977 1218
rect 3880 242 3931 1194
rect 3965 242 3977 1194
rect 3880 218 3977 242
rect 4303 1194 4400 1218
rect 4303 242 4315 1194
rect 4349 242 4400 1194
rect 4303 218 4400 242
rect 4800 1194 4897 1218
rect 4800 242 4851 1194
rect 4885 242 4897 1194
rect 4800 218 4897 242
rect 5223 1194 5320 1218
rect 5223 242 5235 1194
rect 5269 242 5320 1194
rect 5223 218 5320 242
rect 5720 1194 5817 1218
rect 5720 242 5771 1194
rect 5805 242 5817 1194
rect 5720 218 5817 242
rect 6143 1194 6240 1218
rect 6143 242 6155 1194
rect 6189 242 6240 1194
rect 6143 218 6240 242
rect 6640 1194 6737 1218
rect 6640 242 6691 1194
rect 6725 242 6737 1194
rect 6640 218 6737 242
rect -6737 -242 -6640 -218
rect -6737 -1194 -6725 -242
rect -6691 -1194 -6640 -242
rect -6737 -1218 -6640 -1194
rect -6240 -242 -6143 -218
rect -6240 -1194 -6189 -242
rect -6155 -1194 -6143 -242
rect -6240 -1218 -6143 -1194
rect -5817 -242 -5720 -218
rect -5817 -1194 -5805 -242
rect -5771 -1194 -5720 -242
rect -5817 -1218 -5720 -1194
rect -5320 -242 -5223 -218
rect -5320 -1194 -5269 -242
rect -5235 -1194 -5223 -242
rect -5320 -1218 -5223 -1194
rect -4897 -242 -4800 -218
rect -4897 -1194 -4885 -242
rect -4851 -1194 -4800 -242
rect -4897 -1218 -4800 -1194
rect -4400 -242 -4303 -218
rect -4400 -1194 -4349 -242
rect -4315 -1194 -4303 -242
rect -4400 -1218 -4303 -1194
rect -3977 -242 -3880 -218
rect -3977 -1194 -3965 -242
rect -3931 -1194 -3880 -242
rect -3977 -1218 -3880 -1194
rect -3480 -242 -3383 -218
rect -3480 -1194 -3429 -242
rect -3395 -1194 -3383 -242
rect -3480 -1218 -3383 -1194
rect -3057 -242 -2960 -218
rect -3057 -1194 -3045 -242
rect -3011 -1194 -2960 -242
rect -3057 -1218 -2960 -1194
rect -2560 -242 -2463 -218
rect -2560 -1194 -2509 -242
rect -2475 -1194 -2463 -242
rect -2560 -1218 -2463 -1194
rect -2137 -242 -2040 -218
rect -2137 -1194 -2125 -242
rect -2091 -1194 -2040 -242
rect -2137 -1218 -2040 -1194
rect -1640 -242 -1543 -218
rect -1640 -1194 -1589 -242
rect -1555 -1194 -1543 -242
rect -1640 -1218 -1543 -1194
rect -1217 -242 -1120 -218
rect -1217 -1194 -1205 -242
rect -1171 -1194 -1120 -242
rect -1217 -1218 -1120 -1194
rect -720 -242 -623 -218
rect -720 -1194 -669 -242
rect -635 -1194 -623 -242
rect -720 -1218 -623 -1194
rect -297 -242 -200 -218
rect -297 -1194 -285 -242
rect -251 -1194 -200 -242
rect -297 -1218 -200 -1194
rect 200 -242 297 -218
rect 200 -1194 251 -242
rect 285 -1194 297 -242
rect 200 -1218 297 -1194
rect 623 -242 720 -218
rect 623 -1194 635 -242
rect 669 -1194 720 -242
rect 623 -1218 720 -1194
rect 1120 -242 1217 -218
rect 1120 -1194 1171 -242
rect 1205 -1194 1217 -242
rect 1120 -1218 1217 -1194
rect 1543 -242 1640 -218
rect 1543 -1194 1555 -242
rect 1589 -1194 1640 -242
rect 1543 -1218 1640 -1194
rect 2040 -242 2137 -218
rect 2040 -1194 2091 -242
rect 2125 -1194 2137 -242
rect 2040 -1218 2137 -1194
rect 2463 -242 2560 -218
rect 2463 -1194 2475 -242
rect 2509 -1194 2560 -242
rect 2463 -1218 2560 -1194
rect 2960 -242 3057 -218
rect 2960 -1194 3011 -242
rect 3045 -1194 3057 -242
rect 2960 -1218 3057 -1194
rect 3383 -242 3480 -218
rect 3383 -1194 3395 -242
rect 3429 -1194 3480 -242
rect 3383 -1218 3480 -1194
rect 3880 -242 3977 -218
rect 3880 -1194 3931 -242
rect 3965 -1194 3977 -242
rect 3880 -1218 3977 -1194
rect 4303 -242 4400 -218
rect 4303 -1194 4315 -242
rect 4349 -1194 4400 -242
rect 4303 -1218 4400 -1194
rect 4800 -242 4897 -218
rect 4800 -1194 4851 -242
rect 4885 -1194 4897 -242
rect 4800 -1218 4897 -1194
rect 5223 -242 5320 -218
rect 5223 -1194 5235 -242
rect 5269 -1194 5320 -242
rect 5223 -1218 5320 -1194
rect 5720 -242 5817 -218
rect 5720 -1194 5771 -242
rect 5805 -1194 5817 -242
rect 5720 -1218 5817 -1194
rect 6143 -242 6240 -218
rect 6143 -1194 6155 -242
rect 6189 -1194 6240 -242
rect 6143 -1218 6240 -1194
rect 6640 -242 6737 -218
rect 6640 -1194 6691 -242
rect 6725 -1194 6737 -242
rect 6640 -1218 6737 -1194
<< psubdiffcont >>
rect -6751 1349 6751 1383
rect -6847 -1287 -6813 1287
rect 6813 -1287 6847 1287
rect -6751 -1383 6751 -1349
<< nsubdiffcont >>
rect -6725 242 -6691 1194
rect -6189 242 -6155 1194
rect -5805 242 -5771 1194
rect -5269 242 -5235 1194
rect -4885 242 -4851 1194
rect -4349 242 -4315 1194
rect -3965 242 -3931 1194
rect -3429 242 -3395 1194
rect -3045 242 -3011 1194
rect -2509 242 -2475 1194
rect -2125 242 -2091 1194
rect -1589 242 -1555 1194
rect -1205 242 -1171 1194
rect -669 242 -635 1194
rect -285 242 -251 1194
rect 251 242 285 1194
rect 635 242 669 1194
rect 1171 242 1205 1194
rect 1555 242 1589 1194
rect 2091 242 2125 1194
rect 2475 242 2509 1194
rect 3011 242 3045 1194
rect 3395 242 3429 1194
rect 3931 242 3965 1194
rect 4315 242 4349 1194
rect 4851 242 4885 1194
rect 5235 242 5269 1194
rect 5771 242 5805 1194
rect 6155 242 6189 1194
rect 6691 242 6725 1194
rect -6725 -1194 -6691 -242
rect -6189 -1194 -6155 -242
rect -5805 -1194 -5771 -242
rect -5269 -1194 -5235 -242
rect -4885 -1194 -4851 -242
rect -4349 -1194 -4315 -242
rect -3965 -1194 -3931 -242
rect -3429 -1194 -3395 -242
rect -3045 -1194 -3011 -242
rect -2509 -1194 -2475 -242
rect -2125 -1194 -2091 -242
rect -1589 -1194 -1555 -242
rect -1205 -1194 -1171 -242
rect -669 -1194 -635 -242
rect -285 -1194 -251 -242
rect 251 -1194 285 -242
rect 635 -1194 669 -242
rect 1171 -1194 1205 -242
rect 1555 -1194 1589 -242
rect 2091 -1194 2125 -242
rect 2475 -1194 2509 -242
rect 3011 -1194 3045 -242
rect 3395 -1194 3429 -242
rect 3931 -1194 3965 -242
rect 4315 -1194 4349 -242
rect 4851 -1194 4885 -242
rect 5235 -1194 5269 -242
rect 5771 -1194 5805 -242
rect 6155 -1194 6189 -242
rect 6691 -1194 6725 -242
<< poly >>
rect -6640 1290 -6240 1306
rect -6640 1256 -6624 1290
rect -6256 1256 -6240 1290
rect -6640 1218 -6240 1256
rect -5720 1290 -5320 1306
rect -5720 1256 -5704 1290
rect -5336 1256 -5320 1290
rect -5720 1218 -5320 1256
rect -4800 1290 -4400 1306
rect -4800 1256 -4784 1290
rect -4416 1256 -4400 1290
rect -4800 1218 -4400 1256
rect -3880 1290 -3480 1306
rect -3880 1256 -3864 1290
rect -3496 1256 -3480 1290
rect -3880 1218 -3480 1256
rect -2960 1290 -2560 1306
rect -2960 1256 -2944 1290
rect -2576 1256 -2560 1290
rect -2960 1218 -2560 1256
rect -2040 1290 -1640 1306
rect -2040 1256 -2024 1290
rect -1656 1256 -1640 1290
rect -2040 1218 -1640 1256
rect -1120 1290 -720 1306
rect -1120 1256 -1104 1290
rect -736 1256 -720 1290
rect -1120 1218 -720 1256
rect -200 1290 200 1306
rect -200 1256 -184 1290
rect 184 1256 200 1290
rect -200 1218 200 1256
rect 720 1290 1120 1306
rect 720 1256 736 1290
rect 1104 1256 1120 1290
rect 720 1218 1120 1256
rect 1640 1290 2040 1306
rect 1640 1256 1656 1290
rect 2024 1256 2040 1290
rect 1640 1218 2040 1256
rect 2560 1290 2960 1306
rect 2560 1256 2576 1290
rect 2944 1256 2960 1290
rect 2560 1218 2960 1256
rect 3480 1290 3880 1306
rect 3480 1256 3496 1290
rect 3864 1256 3880 1290
rect 3480 1218 3880 1256
rect 4400 1290 4800 1306
rect 4400 1256 4416 1290
rect 4784 1256 4800 1290
rect 4400 1218 4800 1256
rect 5320 1290 5720 1306
rect 5320 1256 5336 1290
rect 5704 1256 5720 1290
rect 5320 1218 5720 1256
rect 6240 1290 6640 1306
rect 6240 1256 6256 1290
rect 6624 1256 6640 1290
rect 6240 1218 6640 1256
rect -6640 180 -6240 218
rect -6640 146 -6624 180
rect -6256 146 -6240 180
rect -6640 130 -6240 146
rect -5720 180 -5320 218
rect -5720 146 -5704 180
rect -5336 146 -5320 180
rect -5720 130 -5320 146
rect -4800 180 -4400 218
rect -4800 146 -4784 180
rect -4416 146 -4400 180
rect -4800 130 -4400 146
rect -3880 180 -3480 218
rect -3880 146 -3864 180
rect -3496 146 -3480 180
rect -3880 130 -3480 146
rect -2960 180 -2560 218
rect -2960 146 -2944 180
rect -2576 146 -2560 180
rect -2960 130 -2560 146
rect -2040 180 -1640 218
rect -2040 146 -2024 180
rect -1656 146 -1640 180
rect -2040 130 -1640 146
rect -1120 180 -720 218
rect -1120 146 -1104 180
rect -736 146 -720 180
rect -1120 130 -720 146
rect -200 180 200 218
rect -200 146 -184 180
rect 184 146 200 180
rect -200 130 200 146
rect 720 180 1120 218
rect 720 146 736 180
rect 1104 146 1120 180
rect 720 130 1120 146
rect 1640 180 2040 218
rect 1640 146 1656 180
rect 2024 146 2040 180
rect 1640 130 2040 146
rect 2560 180 2960 218
rect 2560 146 2576 180
rect 2944 146 2960 180
rect 2560 130 2960 146
rect 3480 180 3880 218
rect 3480 146 3496 180
rect 3864 146 3880 180
rect 3480 130 3880 146
rect 4400 180 4800 218
rect 4400 146 4416 180
rect 4784 146 4800 180
rect 4400 130 4800 146
rect 5320 180 5720 218
rect 5320 146 5336 180
rect 5704 146 5720 180
rect 5320 130 5720 146
rect 6240 180 6640 218
rect 6240 146 6256 180
rect 6624 146 6640 180
rect 6240 130 6640 146
rect -6640 -146 -6240 -130
rect -6640 -180 -6624 -146
rect -6256 -180 -6240 -146
rect -6640 -218 -6240 -180
rect -5720 -146 -5320 -130
rect -5720 -180 -5704 -146
rect -5336 -180 -5320 -146
rect -5720 -218 -5320 -180
rect -4800 -146 -4400 -130
rect -4800 -180 -4784 -146
rect -4416 -180 -4400 -146
rect -4800 -218 -4400 -180
rect -3880 -146 -3480 -130
rect -3880 -180 -3864 -146
rect -3496 -180 -3480 -146
rect -3880 -218 -3480 -180
rect -2960 -146 -2560 -130
rect -2960 -180 -2944 -146
rect -2576 -180 -2560 -146
rect -2960 -218 -2560 -180
rect -2040 -146 -1640 -130
rect -2040 -180 -2024 -146
rect -1656 -180 -1640 -146
rect -2040 -218 -1640 -180
rect -1120 -146 -720 -130
rect -1120 -180 -1104 -146
rect -736 -180 -720 -146
rect -1120 -218 -720 -180
rect -200 -146 200 -130
rect -200 -180 -184 -146
rect 184 -180 200 -146
rect -200 -218 200 -180
rect 720 -146 1120 -130
rect 720 -180 736 -146
rect 1104 -180 1120 -146
rect 720 -218 1120 -180
rect 1640 -146 2040 -130
rect 1640 -180 1656 -146
rect 2024 -180 2040 -146
rect 1640 -218 2040 -180
rect 2560 -146 2960 -130
rect 2560 -180 2576 -146
rect 2944 -180 2960 -146
rect 2560 -218 2960 -180
rect 3480 -146 3880 -130
rect 3480 -180 3496 -146
rect 3864 -180 3880 -146
rect 3480 -218 3880 -180
rect 4400 -146 4800 -130
rect 4400 -180 4416 -146
rect 4784 -180 4800 -146
rect 4400 -218 4800 -180
rect 5320 -146 5720 -130
rect 5320 -180 5336 -146
rect 5704 -180 5720 -146
rect 5320 -218 5720 -180
rect 6240 -146 6640 -130
rect 6240 -180 6256 -146
rect 6624 -180 6640 -146
rect 6240 -218 6640 -180
rect -6640 -1256 -6240 -1218
rect -6640 -1290 -6624 -1256
rect -6256 -1290 -6240 -1256
rect -6640 -1306 -6240 -1290
rect -5720 -1256 -5320 -1218
rect -5720 -1290 -5704 -1256
rect -5336 -1290 -5320 -1256
rect -5720 -1306 -5320 -1290
rect -4800 -1256 -4400 -1218
rect -4800 -1290 -4784 -1256
rect -4416 -1290 -4400 -1256
rect -4800 -1306 -4400 -1290
rect -3880 -1256 -3480 -1218
rect -3880 -1290 -3864 -1256
rect -3496 -1290 -3480 -1256
rect -3880 -1306 -3480 -1290
rect -2960 -1256 -2560 -1218
rect -2960 -1290 -2944 -1256
rect -2576 -1290 -2560 -1256
rect -2960 -1306 -2560 -1290
rect -2040 -1256 -1640 -1218
rect -2040 -1290 -2024 -1256
rect -1656 -1290 -1640 -1256
rect -2040 -1306 -1640 -1290
rect -1120 -1256 -720 -1218
rect -1120 -1290 -1104 -1256
rect -736 -1290 -720 -1256
rect -1120 -1306 -720 -1290
rect -200 -1256 200 -1218
rect -200 -1290 -184 -1256
rect 184 -1290 200 -1256
rect -200 -1306 200 -1290
rect 720 -1256 1120 -1218
rect 720 -1290 736 -1256
rect 1104 -1290 1120 -1256
rect 720 -1306 1120 -1290
rect 1640 -1256 2040 -1218
rect 1640 -1290 1656 -1256
rect 2024 -1290 2040 -1256
rect 1640 -1306 2040 -1290
rect 2560 -1256 2960 -1218
rect 2560 -1290 2576 -1256
rect 2944 -1290 2960 -1256
rect 2560 -1306 2960 -1290
rect 3480 -1256 3880 -1218
rect 3480 -1290 3496 -1256
rect 3864 -1290 3880 -1256
rect 3480 -1306 3880 -1290
rect 4400 -1256 4800 -1218
rect 4400 -1290 4416 -1256
rect 4784 -1290 4800 -1256
rect 4400 -1306 4800 -1290
rect 5320 -1256 5720 -1218
rect 5320 -1290 5336 -1256
rect 5704 -1290 5720 -1256
rect 5320 -1306 5720 -1290
rect 6240 -1256 6640 -1218
rect 6240 -1290 6256 -1256
rect 6624 -1290 6640 -1256
rect 6240 -1306 6640 -1290
<< polycont >>
rect -6624 1256 -6256 1290
rect -5704 1256 -5336 1290
rect -4784 1256 -4416 1290
rect -3864 1256 -3496 1290
rect -2944 1256 -2576 1290
rect -2024 1256 -1656 1290
rect -1104 1256 -736 1290
rect -184 1256 184 1290
rect 736 1256 1104 1290
rect 1656 1256 2024 1290
rect 2576 1256 2944 1290
rect 3496 1256 3864 1290
rect 4416 1256 4784 1290
rect 5336 1256 5704 1290
rect 6256 1256 6624 1290
rect -6624 146 -6256 180
rect -5704 146 -5336 180
rect -4784 146 -4416 180
rect -3864 146 -3496 180
rect -2944 146 -2576 180
rect -2024 146 -1656 180
rect -1104 146 -736 180
rect -184 146 184 180
rect 736 146 1104 180
rect 1656 146 2024 180
rect 2576 146 2944 180
rect 3496 146 3864 180
rect 4416 146 4784 180
rect 5336 146 5704 180
rect 6256 146 6624 180
rect -6624 -180 -6256 -146
rect -5704 -180 -5336 -146
rect -4784 -180 -4416 -146
rect -3864 -180 -3496 -146
rect -2944 -180 -2576 -146
rect -2024 -180 -1656 -146
rect -1104 -180 -736 -146
rect -184 -180 184 -146
rect 736 -180 1104 -146
rect 1656 -180 2024 -146
rect 2576 -180 2944 -146
rect 3496 -180 3864 -146
rect 4416 -180 4784 -146
rect 5336 -180 5704 -146
rect 6256 -180 6624 -146
rect -6624 -1290 -6256 -1256
rect -5704 -1290 -5336 -1256
rect -4784 -1290 -4416 -1256
rect -3864 -1290 -3496 -1256
rect -2944 -1290 -2576 -1256
rect -2024 -1290 -1656 -1256
rect -1104 -1290 -736 -1256
rect -184 -1290 184 -1256
rect 736 -1290 1104 -1256
rect 1656 -1290 2024 -1256
rect 2576 -1290 2944 -1256
rect 3496 -1290 3864 -1256
rect 4416 -1290 4784 -1256
rect 5336 -1290 5704 -1256
rect 6256 -1290 6624 -1256
<< locali >>
rect -6847 1349 -6751 1383
rect 6751 1349 6847 1383
rect -6847 1287 -6813 1349
rect -6640 1256 -6624 1290
rect -6256 1256 -6240 1290
rect -5720 1256 -5704 1290
rect -5336 1256 -5320 1290
rect -4800 1256 -4784 1290
rect -4416 1256 -4400 1290
rect -3880 1256 -3864 1290
rect -3496 1256 -3480 1290
rect -2960 1256 -2944 1290
rect -2576 1256 -2560 1290
rect -2040 1256 -2024 1290
rect -1656 1256 -1640 1290
rect -1120 1256 -1104 1290
rect -736 1256 -720 1290
rect -200 1256 -184 1290
rect 184 1256 200 1290
rect 720 1256 736 1290
rect 1104 1256 1120 1290
rect 1640 1256 1656 1290
rect 2024 1256 2040 1290
rect 2560 1256 2576 1290
rect 2944 1256 2960 1290
rect 3480 1256 3496 1290
rect 3864 1256 3880 1290
rect 4400 1256 4416 1290
rect 4784 1256 4800 1290
rect 5320 1256 5336 1290
rect 5704 1256 5720 1290
rect 6240 1256 6256 1290
rect 6624 1256 6640 1290
rect 6813 1287 6847 1349
rect -6725 1194 -6691 1210
rect -6725 226 -6691 242
rect -6189 1194 -6155 1210
rect -6189 226 -6155 242
rect -5805 1194 -5771 1210
rect -5805 226 -5771 242
rect -5269 1194 -5235 1210
rect -5269 226 -5235 242
rect -4885 1194 -4851 1210
rect -4885 226 -4851 242
rect -4349 1194 -4315 1210
rect -4349 226 -4315 242
rect -3965 1194 -3931 1210
rect -3965 226 -3931 242
rect -3429 1194 -3395 1210
rect -3429 226 -3395 242
rect -3045 1194 -3011 1210
rect -3045 226 -3011 242
rect -2509 1194 -2475 1210
rect -2509 226 -2475 242
rect -2125 1194 -2091 1210
rect -2125 226 -2091 242
rect -1589 1194 -1555 1210
rect -1589 226 -1555 242
rect -1205 1194 -1171 1210
rect -1205 226 -1171 242
rect -669 1194 -635 1210
rect -669 226 -635 242
rect -285 1194 -251 1210
rect -285 226 -251 242
rect 251 1194 285 1210
rect 251 226 285 242
rect 635 1194 669 1210
rect 635 226 669 242
rect 1171 1194 1205 1210
rect 1171 226 1205 242
rect 1555 1194 1589 1210
rect 1555 226 1589 242
rect 2091 1194 2125 1210
rect 2091 226 2125 242
rect 2475 1194 2509 1210
rect 2475 226 2509 242
rect 3011 1194 3045 1210
rect 3011 226 3045 242
rect 3395 1194 3429 1210
rect 3395 226 3429 242
rect 3931 1194 3965 1210
rect 3931 226 3965 242
rect 4315 1194 4349 1210
rect 4315 226 4349 242
rect 4851 1194 4885 1210
rect 4851 226 4885 242
rect 5235 1194 5269 1210
rect 5235 226 5269 242
rect 5771 1194 5805 1210
rect 5771 226 5805 242
rect 6155 1194 6189 1210
rect 6155 226 6189 242
rect 6691 1194 6725 1210
rect 6691 226 6725 242
rect -6640 146 -6624 180
rect -6256 146 -6240 180
rect -5720 146 -5704 180
rect -5336 146 -5320 180
rect -4800 146 -4784 180
rect -4416 146 -4400 180
rect -3880 146 -3864 180
rect -3496 146 -3480 180
rect -2960 146 -2944 180
rect -2576 146 -2560 180
rect -2040 146 -2024 180
rect -1656 146 -1640 180
rect -1120 146 -1104 180
rect -736 146 -720 180
rect -200 146 -184 180
rect 184 146 200 180
rect 720 146 736 180
rect 1104 146 1120 180
rect 1640 146 1656 180
rect 2024 146 2040 180
rect 2560 146 2576 180
rect 2944 146 2960 180
rect 3480 146 3496 180
rect 3864 146 3880 180
rect 4400 146 4416 180
rect 4784 146 4800 180
rect 5320 146 5336 180
rect 5704 146 5720 180
rect 6240 146 6256 180
rect 6624 146 6640 180
rect -6640 -180 -6624 -146
rect -6256 -180 -6240 -146
rect -5720 -180 -5704 -146
rect -5336 -180 -5320 -146
rect -4800 -180 -4784 -146
rect -4416 -180 -4400 -146
rect -3880 -180 -3864 -146
rect -3496 -180 -3480 -146
rect -2960 -180 -2944 -146
rect -2576 -180 -2560 -146
rect -2040 -180 -2024 -146
rect -1656 -180 -1640 -146
rect -1120 -180 -1104 -146
rect -736 -180 -720 -146
rect -200 -180 -184 -146
rect 184 -180 200 -146
rect 720 -180 736 -146
rect 1104 -180 1120 -146
rect 1640 -180 1656 -146
rect 2024 -180 2040 -146
rect 2560 -180 2576 -146
rect 2944 -180 2960 -146
rect 3480 -180 3496 -146
rect 3864 -180 3880 -146
rect 4400 -180 4416 -146
rect 4784 -180 4800 -146
rect 5320 -180 5336 -146
rect 5704 -180 5720 -146
rect 6240 -180 6256 -146
rect 6624 -180 6640 -146
rect -6725 -242 -6691 -226
rect -6725 -1210 -6691 -1194
rect -6189 -242 -6155 -226
rect -6189 -1210 -6155 -1194
rect -5805 -242 -5771 -226
rect -5805 -1210 -5771 -1194
rect -5269 -242 -5235 -226
rect -5269 -1210 -5235 -1194
rect -4885 -242 -4851 -226
rect -4885 -1210 -4851 -1194
rect -4349 -242 -4315 -226
rect -4349 -1210 -4315 -1194
rect -3965 -242 -3931 -226
rect -3965 -1210 -3931 -1194
rect -3429 -242 -3395 -226
rect -3429 -1210 -3395 -1194
rect -3045 -242 -3011 -226
rect -3045 -1210 -3011 -1194
rect -2509 -242 -2475 -226
rect -2509 -1210 -2475 -1194
rect -2125 -242 -2091 -226
rect -2125 -1210 -2091 -1194
rect -1589 -242 -1555 -226
rect -1589 -1210 -1555 -1194
rect -1205 -242 -1171 -226
rect -1205 -1210 -1171 -1194
rect -669 -242 -635 -226
rect -669 -1210 -635 -1194
rect -285 -242 -251 -226
rect -285 -1210 -251 -1194
rect 251 -242 285 -226
rect 251 -1210 285 -1194
rect 635 -242 669 -226
rect 635 -1210 669 -1194
rect 1171 -242 1205 -226
rect 1171 -1210 1205 -1194
rect 1555 -242 1589 -226
rect 1555 -1210 1589 -1194
rect 2091 -242 2125 -226
rect 2091 -1210 2125 -1194
rect 2475 -242 2509 -226
rect 2475 -1210 2509 -1194
rect 3011 -242 3045 -226
rect 3011 -1210 3045 -1194
rect 3395 -242 3429 -226
rect 3395 -1210 3429 -1194
rect 3931 -242 3965 -226
rect 3931 -1210 3965 -1194
rect 4315 -242 4349 -226
rect 4315 -1210 4349 -1194
rect 4851 -242 4885 -226
rect 4851 -1210 4885 -1194
rect 5235 -242 5269 -226
rect 5235 -1210 5269 -1194
rect 5771 -242 5805 -226
rect 5771 -1210 5805 -1194
rect 6155 -242 6189 -226
rect 6155 -1210 6189 -1194
rect 6691 -242 6725 -226
rect 6691 -1210 6725 -1194
rect -6847 -1349 -6813 -1287
rect -6640 -1290 -6624 -1256
rect -6256 -1290 -6240 -1256
rect -5720 -1290 -5704 -1256
rect -5336 -1290 -5320 -1256
rect -4800 -1290 -4784 -1256
rect -4416 -1290 -4400 -1256
rect -3880 -1290 -3864 -1256
rect -3496 -1290 -3480 -1256
rect -2960 -1290 -2944 -1256
rect -2576 -1290 -2560 -1256
rect -2040 -1290 -2024 -1256
rect -1656 -1290 -1640 -1256
rect -1120 -1290 -1104 -1256
rect -736 -1290 -720 -1256
rect -200 -1290 -184 -1256
rect 184 -1290 200 -1256
rect 720 -1290 736 -1256
rect 1104 -1290 1120 -1256
rect 1640 -1290 1656 -1256
rect 2024 -1290 2040 -1256
rect 2560 -1290 2576 -1256
rect 2944 -1290 2960 -1256
rect 3480 -1290 3496 -1256
rect 3864 -1290 3880 -1256
rect 4400 -1290 4416 -1256
rect 4784 -1290 4800 -1256
rect 5320 -1290 5336 -1256
rect 5704 -1290 5720 -1256
rect 6240 -1290 6256 -1256
rect 6624 -1290 6640 -1256
rect 6813 -1349 6847 -1287
rect -6847 -1383 -6751 -1349
rect 6751 -1383 6847 -1349
<< viali >>
rect -6624 1256 -6256 1290
rect -5704 1256 -5336 1290
rect -4784 1256 -4416 1290
rect -3864 1256 -3496 1290
rect -2944 1256 -2576 1290
rect -2024 1256 -1656 1290
rect -1104 1256 -736 1290
rect -184 1256 184 1290
rect 736 1256 1104 1290
rect 1656 1256 2024 1290
rect 2576 1256 2944 1290
rect 3496 1256 3864 1290
rect 4416 1256 4784 1290
rect 5336 1256 5704 1290
rect 6256 1256 6624 1290
rect -6725 242 -6691 1194
rect -6189 242 -6155 1194
rect -5805 242 -5771 1194
rect -5269 242 -5235 1194
rect -4885 242 -4851 1194
rect -4349 242 -4315 1194
rect -3965 242 -3931 1194
rect -3429 242 -3395 1194
rect -3045 242 -3011 1194
rect -2509 242 -2475 1194
rect -2125 242 -2091 1194
rect -1589 242 -1555 1194
rect -1205 242 -1171 1194
rect -669 242 -635 1194
rect -285 242 -251 1194
rect 251 242 285 1194
rect 635 242 669 1194
rect 1171 242 1205 1194
rect 1555 242 1589 1194
rect 2091 242 2125 1194
rect 2475 242 2509 1194
rect 3011 242 3045 1194
rect 3395 242 3429 1194
rect 3931 242 3965 1194
rect 4315 242 4349 1194
rect 4851 242 4885 1194
rect 5235 242 5269 1194
rect 5771 242 5805 1194
rect 6155 242 6189 1194
rect 6691 242 6725 1194
rect -6624 146 -6256 180
rect -5704 146 -5336 180
rect -4784 146 -4416 180
rect -3864 146 -3496 180
rect -2944 146 -2576 180
rect -2024 146 -1656 180
rect -1104 146 -736 180
rect -184 146 184 180
rect 736 146 1104 180
rect 1656 146 2024 180
rect 2576 146 2944 180
rect 3496 146 3864 180
rect 4416 146 4784 180
rect 5336 146 5704 180
rect 6256 146 6624 180
rect -6624 -180 -6256 -146
rect -5704 -180 -5336 -146
rect -4784 -180 -4416 -146
rect -3864 -180 -3496 -146
rect -2944 -180 -2576 -146
rect -2024 -180 -1656 -146
rect -1104 -180 -736 -146
rect -184 -180 184 -146
rect 736 -180 1104 -146
rect 1656 -180 2024 -146
rect 2576 -180 2944 -146
rect 3496 -180 3864 -146
rect 4416 -180 4784 -146
rect 5336 -180 5704 -146
rect 6256 -180 6624 -146
rect -6725 -1194 -6691 -242
rect -6189 -1194 -6155 -242
rect -5805 -1194 -5771 -242
rect -5269 -1194 -5235 -242
rect -4885 -1194 -4851 -242
rect -4349 -1194 -4315 -242
rect -3965 -1194 -3931 -242
rect -3429 -1194 -3395 -242
rect -3045 -1194 -3011 -242
rect -2509 -1194 -2475 -242
rect -2125 -1194 -2091 -242
rect -1589 -1194 -1555 -242
rect -1205 -1194 -1171 -242
rect -669 -1194 -635 -242
rect -285 -1194 -251 -242
rect 251 -1194 285 -242
rect 635 -1194 669 -242
rect 1171 -1194 1205 -242
rect 1555 -1194 1589 -242
rect 2091 -1194 2125 -242
rect 2475 -1194 2509 -242
rect 3011 -1194 3045 -242
rect 3395 -1194 3429 -242
rect 3931 -1194 3965 -242
rect 4315 -1194 4349 -242
rect 4851 -1194 4885 -242
rect 5235 -1194 5269 -242
rect 5771 -1194 5805 -242
rect 6155 -1194 6189 -242
rect 6691 -1194 6725 -242
rect -6624 -1290 -6256 -1256
rect -5704 -1290 -5336 -1256
rect -4784 -1290 -4416 -1256
rect -3864 -1290 -3496 -1256
rect -2944 -1290 -2576 -1256
rect -2024 -1290 -1656 -1256
rect -1104 -1290 -736 -1256
rect -184 -1290 184 -1256
rect 736 -1290 1104 -1256
rect 1656 -1290 2024 -1256
rect 2576 -1290 2944 -1256
rect 3496 -1290 3864 -1256
rect 4416 -1290 4784 -1256
rect 5336 -1290 5704 -1256
rect 6256 -1290 6624 -1256
<< metal1 >>
rect -6636 1290 -6244 1296
rect -6636 1256 -6624 1290
rect -6256 1256 -6244 1290
rect -6636 1250 -6244 1256
rect -5716 1290 -5324 1296
rect -5716 1256 -5704 1290
rect -5336 1256 -5324 1290
rect -5716 1250 -5324 1256
rect -4796 1290 -4404 1296
rect -4796 1256 -4784 1290
rect -4416 1256 -4404 1290
rect -4796 1250 -4404 1256
rect -3876 1290 -3484 1296
rect -3876 1256 -3864 1290
rect -3496 1256 -3484 1290
rect -3876 1250 -3484 1256
rect -2956 1290 -2564 1296
rect -2956 1256 -2944 1290
rect -2576 1256 -2564 1290
rect -2956 1250 -2564 1256
rect -2036 1290 -1644 1296
rect -2036 1256 -2024 1290
rect -1656 1256 -1644 1290
rect -2036 1250 -1644 1256
rect -1116 1290 -724 1296
rect -1116 1256 -1104 1290
rect -736 1256 -724 1290
rect -1116 1250 -724 1256
rect -196 1290 196 1296
rect -196 1256 -184 1290
rect 184 1256 196 1290
rect -196 1250 196 1256
rect 724 1290 1116 1296
rect 724 1256 736 1290
rect 1104 1256 1116 1290
rect 724 1250 1116 1256
rect 1644 1290 2036 1296
rect 1644 1256 1656 1290
rect 2024 1256 2036 1290
rect 1644 1250 2036 1256
rect 2564 1290 2956 1296
rect 2564 1256 2576 1290
rect 2944 1256 2956 1290
rect 2564 1250 2956 1256
rect 3484 1290 3876 1296
rect 3484 1256 3496 1290
rect 3864 1256 3876 1290
rect 3484 1250 3876 1256
rect 4404 1290 4796 1296
rect 4404 1256 4416 1290
rect 4784 1256 4796 1290
rect 4404 1250 4796 1256
rect 5324 1290 5716 1296
rect 5324 1256 5336 1290
rect 5704 1256 5716 1290
rect 5324 1250 5716 1256
rect 6244 1290 6636 1296
rect 6244 1256 6256 1290
rect 6624 1256 6636 1290
rect 6244 1250 6636 1256
rect -6731 1194 -6685 1206
rect -6731 242 -6725 1194
rect -6691 242 -6685 1194
rect -6731 230 -6685 242
rect -6195 1194 -6149 1206
rect -6195 242 -6189 1194
rect -6155 242 -6149 1194
rect -6195 230 -6149 242
rect -5811 1194 -5765 1206
rect -5811 242 -5805 1194
rect -5771 242 -5765 1194
rect -5811 230 -5765 242
rect -5275 1194 -5229 1206
rect -5275 242 -5269 1194
rect -5235 242 -5229 1194
rect -5275 230 -5229 242
rect -4891 1194 -4845 1206
rect -4891 242 -4885 1194
rect -4851 242 -4845 1194
rect -4891 230 -4845 242
rect -4355 1194 -4309 1206
rect -4355 242 -4349 1194
rect -4315 242 -4309 1194
rect -4355 230 -4309 242
rect -3971 1194 -3925 1206
rect -3971 242 -3965 1194
rect -3931 242 -3925 1194
rect -3971 230 -3925 242
rect -3435 1194 -3389 1206
rect -3435 242 -3429 1194
rect -3395 242 -3389 1194
rect -3435 230 -3389 242
rect -3051 1194 -3005 1206
rect -3051 242 -3045 1194
rect -3011 242 -3005 1194
rect -3051 230 -3005 242
rect -2515 1194 -2469 1206
rect -2515 242 -2509 1194
rect -2475 242 -2469 1194
rect -2515 230 -2469 242
rect -2131 1194 -2085 1206
rect -2131 242 -2125 1194
rect -2091 242 -2085 1194
rect -2131 230 -2085 242
rect -1595 1194 -1549 1206
rect -1595 242 -1589 1194
rect -1555 242 -1549 1194
rect -1595 230 -1549 242
rect -1211 1194 -1165 1206
rect -1211 242 -1205 1194
rect -1171 242 -1165 1194
rect -1211 230 -1165 242
rect -675 1194 -629 1206
rect -675 242 -669 1194
rect -635 242 -629 1194
rect -675 230 -629 242
rect -291 1194 -245 1206
rect -291 242 -285 1194
rect -251 242 -245 1194
rect -291 230 -245 242
rect 245 1194 291 1206
rect 245 242 251 1194
rect 285 242 291 1194
rect 245 230 291 242
rect 629 1194 675 1206
rect 629 242 635 1194
rect 669 242 675 1194
rect 629 230 675 242
rect 1165 1194 1211 1206
rect 1165 242 1171 1194
rect 1205 242 1211 1194
rect 1165 230 1211 242
rect 1549 1194 1595 1206
rect 1549 242 1555 1194
rect 1589 242 1595 1194
rect 1549 230 1595 242
rect 2085 1194 2131 1206
rect 2085 242 2091 1194
rect 2125 242 2131 1194
rect 2085 230 2131 242
rect 2469 1194 2515 1206
rect 2469 242 2475 1194
rect 2509 242 2515 1194
rect 2469 230 2515 242
rect 3005 1194 3051 1206
rect 3005 242 3011 1194
rect 3045 242 3051 1194
rect 3005 230 3051 242
rect 3389 1194 3435 1206
rect 3389 242 3395 1194
rect 3429 242 3435 1194
rect 3389 230 3435 242
rect 3925 1194 3971 1206
rect 3925 242 3931 1194
rect 3965 242 3971 1194
rect 3925 230 3971 242
rect 4309 1194 4355 1206
rect 4309 242 4315 1194
rect 4349 242 4355 1194
rect 4309 230 4355 242
rect 4845 1194 4891 1206
rect 4845 242 4851 1194
rect 4885 242 4891 1194
rect 4845 230 4891 242
rect 5229 1194 5275 1206
rect 5229 242 5235 1194
rect 5269 242 5275 1194
rect 5229 230 5275 242
rect 5765 1194 5811 1206
rect 5765 242 5771 1194
rect 5805 242 5811 1194
rect 5765 230 5811 242
rect 6149 1194 6195 1206
rect 6149 242 6155 1194
rect 6189 242 6195 1194
rect 6149 230 6195 242
rect 6685 1194 6731 1206
rect 6685 242 6691 1194
rect 6725 242 6731 1194
rect 6685 230 6731 242
rect -6636 180 -6244 186
rect -6636 146 -6624 180
rect -6256 146 -6244 180
rect -6636 140 -6244 146
rect -5716 180 -5324 186
rect -5716 146 -5704 180
rect -5336 146 -5324 180
rect -5716 140 -5324 146
rect -4796 180 -4404 186
rect -4796 146 -4784 180
rect -4416 146 -4404 180
rect -4796 140 -4404 146
rect -3876 180 -3484 186
rect -3876 146 -3864 180
rect -3496 146 -3484 180
rect -3876 140 -3484 146
rect -2956 180 -2564 186
rect -2956 146 -2944 180
rect -2576 146 -2564 180
rect -2956 140 -2564 146
rect -2036 180 -1644 186
rect -2036 146 -2024 180
rect -1656 146 -1644 180
rect -2036 140 -1644 146
rect -1116 180 -724 186
rect -1116 146 -1104 180
rect -736 146 -724 180
rect -1116 140 -724 146
rect -196 180 196 186
rect -196 146 -184 180
rect 184 146 196 180
rect -196 140 196 146
rect 724 180 1116 186
rect 724 146 736 180
rect 1104 146 1116 180
rect 724 140 1116 146
rect 1644 180 2036 186
rect 1644 146 1656 180
rect 2024 146 2036 180
rect 1644 140 2036 146
rect 2564 180 2956 186
rect 2564 146 2576 180
rect 2944 146 2956 180
rect 2564 140 2956 146
rect 3484 180 3876 186
rect 3484 146 3496 180
rect 3864 146 3876 180
rect 3484 140 3876 146
rect 4404 180 4796 186
rect 4404 146 4416 180
rect 4784 146 4796 180
rect 4404 140 4796 146
rect 5324 180 5716 186
rect 5324 146 5336 180
rect 5704 146 5716 180
rect 5324 140 5716 146
rect 6244 180 6636 186
rect 6244 146 6256 180
rect 6624 146 6636 180
rect 6244 140 6636 146
rect -6636 -146 -6244 -140
rect -6636 -180 -6624 -146
rect -6256 -180 -6244 -146
rect -6636 -186 -6244 -180
rect -5716 -146 -5324 -140
rect -5716 -180 -5704 -146
rect -5336 -180 -5324 -146
rect -5716 -186 -5324 -180
rect -4796 -146 -4404 -140
rect -4796 -180 -4784 -146
rect -4416 -180 -4404 -146
rect -4796 -186 -4404 -180
rect -3876 -146 -3484 -140
rect -3876 -180 -3864 -146
rect -3496 -180 -3484 -146
rect -3876 -186 -3484 -180
rect -2956 -146 -2564 -140
rect -2956 -180 -2944 -146
rect -2576 -180 -2564 -146
rect -2956 -186 -2564 -180
rect -2036 -146 -1644 -140
rect -2036 -180 -2024 -146
rect -1656 -180 -1644 -146
rect -2036 -186 -1644 -180
rect -1116 -146 -724 -140
rect -1116 -180 -1104 -146
rect -736 -180 -724 -146
rect -1116 -186 -724 -180
rect -196 -146 196 -140
rect -196 -180 -184 -146
rect 184 -180 196 -146
rect -196 -186 196 -180
rect 724 -146 1116 -140
rect 724 -180 736 -146
rect 1104 -180 1116 -146
rect 724 -186 1116 -180
rect 1644 -146 2036 -140
rect 1644 -180 1656 -146
rect 2024 -180 2036 -146
rect 1644 -186 2036 -180
rect 2564 -146 2956 -140
rect 2564 -180 2576 -146
rect 2944 -180 2956 -146
rect 2564 -186 2956 -180
rect 3484 -146 3876 -140
rect 3484 -180 3496 -146
rect 3864 -180 3876 -146
rect 3484 -186 3876 -180
rect 4404 -146 4796 -140
rect 4404 -180 4416 -146
rect 4784 -180 4796 -146
rect 4404 -186 4796 -180
rect 5324 -146 5716 -140
rect 5324 -180 5336 -146
rect 5704 -180 5716 -146
rect 5324 -186 5716 -180
rect 6244 -146 6636 -140
rect 6244 -180 6256 -146
rect 6624 -180 6636 -146
rect 6244 -186 6636 -180
rect -6731 -242 -6685 -230
rect -6731 -1194 -6725 -242
rect -6691 -1194 -6685 -242
rect -6731 -1206 -6685 -1194
rect -6195 -242 -6149 -230
rect -6195 -1194 -6189 -242
rect -6155 -1194 -6149 -242
rect -6195 -1206 -6149 -1194
rect -5811 -242 -5765 -230
rect -5811 -1194 -5805 -242
rect -5771 -1194 -5765 -242
rect -5811 -1206 -5765 -1194
rect -5275 -242 -5229 -230
rect -5275 -1194 -5269 -242
rect -5235 -1194 -5229 -242
rect -5275 -1206 -5229 -1194
rect -4891 -242 -4845 -230
rect -4891 -1194 -4885 -242
rect -4851 -1194 -4845 -242
rect -4891 -1206 -4845 -1194
rect -4355 -242 -4309 -230
rect -4355 -1194 -4349 -242
rect -4315 -1194 -4309 -242
rect -4355 -1206 -4309 -1194
rect -3971 -242 -3925 -230
rect -3971 -1194 -3965 -242
rect -3931 -1194 -3925 -242
rect -3971 -1206 -3925 -1194
rect -3435 -242 -3389 -230
rect -3435 -1194 -3429 -242
rect -3395 -1194 -3389 -242
rect -3435 -1206 -3389 -1194
rect -3051 -242 -3005 -230
rect -3051 -1194 -3045 -242
rect -3011 -1194 -3005 -242
rect -3051 -1206 -3005 -1194
rect -2515 -242 -2469 -230
rect -2515 -1194 -2509 -242
rect -2475 -1194 -2469 -242
rect -2515 -1206 -2469 -1194
rect -2131 -242 -2085 -230
rect -2131 -1194 -2125 -242
rect -2091 -1194 -2085 -242
rect -2131 -1206 -2085 -1194
rect -1595 -242 -1549 -230
rect -1595 -1194 -1589 -242
rect -1555 -1194 -1549 -242
rect -1595 -1206 -1549 -1194
rect -1211 -242 -1165 -230
rect -1211 -1194 -1205 -242
rect -1171 -1194 -1165 -242
rect -1211 -1206 -1165 -1194
rect -675 -242 -629 -230
rect -675 -1194 -669 -242
rect -635 -1194 -629 -242
rect -675 -1206 -629 -1194
rect -291 -242 -245 -230
rect -291 -1194 -285 -242
rect -251 -1194 -245 -242
rect -291 -1206 -245 -1194
rect 245 -242 291 -230
rect 245 -1194 251 -242
rect 285 -1194 291 -242
rect 245 -1206 291 -1194
rect 629 -242 675 -230
rect 629 -1194 635 -242
rect 669 -1194 675 -242
rect 629 -1206 675 -1194
rect 1165 -242 1211 -230
rect 1165 -1194 1171 -242
rect 1205 -1194 1211 -242
rect 1165 -1206 1211 -1194
rect 1549 -242 1595 -230
rect 1549 -1194 1555 -242
rect 1589 -1194 1595 -242
rect 1549 -1206 1595 -1194
rect 2085 -242 2131 -230
rect 2085 -1194 2091 -242
rect 2125 -1194 2131 -242
rect 2085 -1206 2131 -1194
rect 2469 -242 2515 -230
rect 2469 -1194 2475 -242
rect 2509 -1194 2515 -242
rect 2469 -1206 2515 -1194
rect 3005 -242 3051 -230
rect 3005 -1194 3011 -242
rect 3045 -1194 3051 -242
rect 3005 -1206 3051 -1194
rect 3389 -242 3435 -230
rect 3389 -1194 3395 -242
rect 3429 -1194 3435 -242
rect 3389 -1206 3435 -1194
rect 3925 -242 3971 -230
rect 3925 -1194 3931 -242
rect 3965 -1194 3971 -242
rect 3925 -1206 3971 -1194
rect 4309 -242 4355 -230
rect 4309 -1194 4315 -242
rect 4349 -1194 4355 -242
rect 4309 -1206 4355 -1194
rect 4845 -242 4891 -230
rect 4845 -1194 4851 -242
rect 4885 -1194 4891 -242
rect 4845 -1206 4891 -1194
rect 5229 -242 5275 -230
rect 5229 -1194 5235 -242
rect 5269 -1194 5275 -242
rect 5229 -1206 5275 -1194
rect 5765 -242 5811 -230
rect 5765 -1194 5771 -242
rect 5805 -1194 5811 -242
rect 5765 -1206 5811 -1194
rect 6149 -242 6195 -230
rect 6149 -1194 6155 -242
rect 6189 -1194 6195 -242
rect 6149 -1206 6195 -1194
rect 6685 -242 6731 -230
rect 6685 -1194 6691 -242
rect 6725 -1194 6731 -242
rect 6685 -1206 6731 -1194
rect -6636 -1256 -6244 -1250
rect -6636 -1290 -6624 -1256
rect -6256 -1290 -6244 -1256
rect -6636 -1296 -6244 -1290
rect -5716 -1256 -5324 -1250
rect -5716 -1290 -5704 -1256
rect -5336 -1290 -5324 -1256
rect -5716 -1296 -5324 -1290
rect -4796 -1256 -4404 -1250
rect -4796 -1290 -4784 -1256
rect -4416 -1290 -4404 -1256
rect -4796 -1296 -4404 -1290
rect -3876 -1256 -3484 -1250
rect -3876 -1290 -3864 -1256
rect -3496 -1290 -3484 -1256
rect -3876 -1296 -3484 -1290
rect -2956 -1256 -2564 -1250
rect -2956 -1290 -2944 -1256
rect -2576 -1290 -2564 -1256
rect -2956 -1296 -2564 -1290
rect -2036 -1256 -1644 -1250
rect -2036 -1290 -2024 -1256
rect -1656 -1290 -1644 -1256
rect -2036 -1296 -1644 -1290
rect -1116 -1256 -724 -1250
rect -1116 -1290 -1104 -1256
rect -736 -1290 -724 -1256
rect -1116 -1296 -724 -1290
rect -196 -1256 196 -1250
rect -196 -1290 -184 -1256
rect 184 -1290 196 -1256
rect -196 -1296 196 -1290
rect 724 -1256 1116 -1250
rect 724 -1290 736 -1256
rect 1104 -1290 1116 -1256
rect 724 -1296 1116 -1290
rect 1644 -1256 2036 -1250
rect 1644 -1290 1656 -1256
rect 2024 -1290 2036 -1256
rect 1644 -1296 2036 -1290
rect 2564 -1256 2956 -1250
rect 2564 -1290 2576 -1256
rect 2944 -1290 2956 -1256
rect 2564 -1296 2956 -1290
rect 3484 -1256 3876 -1250
rect 3484 -1290 3496 -1256
rect 3864 -1290 3876 -1256
rect 3484 -1296 3876 -1290
rect 4404 -1256 4796 -1250
rect 4404 -1290 4416 -1256
rect 4784 -1290 4796 -1256
rect 4404 -1296 4796 -1290
rect 5324 -1256 5716 -1250
rect 5324 -1290 5336 -1256
rect 5704 -1290 5716 -1256
rect 5324 -1296 5716 -1290
rect 6244 -1256 6636 -1250
rect 6244 -1290 6256 -1256
rect 6624 -1290 6636 -1256
rect 6244 -1296 6636 -1290
<< properties >>
string FIXED_BBOX -6830 -1366 6830 1366
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 5 l 2 m 2 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
