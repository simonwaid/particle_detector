magic
tech sky130A
magscale 1 2
timestamp 1654771420
<< metal1 >>
rect 51790 18560 51800 18660
rect 51980 18560 51990 18660
rect 52050 18560 52060 18660
rect 52240 18560 52250 18660
rect 49550 14950 49610 14980
rect 92320 9450 92330 9590
rect 92530 9480 92850 9590
rect 92530 9450 92540 9480
rect 49680 8778 49690 9000
rect 49958 8778 49968 9000
rect 67580 3840 67590 4000
rect 67740 3840 67750 4000
<< via1 >>
rect 51800 18560 51980 18660
rect 52060 18560 52240 18660
rect 92330 9450 92530 9590
rect 49690 8778 49958 9000
rect 67590 3840 67740 4000
<< metal2 >>
rect 51800 18660 51980 18670
rect 51800 18550 51980 18560
rect 52060 18660 52240 18670
rect 52060 18550 52240 18560
rect 62300 18150 63700 18560
rect 26770 16240 42160 16380
rect 26770 4130 26910 16240
rect 41840 14240 42160 16240
rect 48810 15130 50480 15320
rect 48820 14240 49020 15130
rect 41840 14050 49020 14240
rect 42040 14040 49020 14050
rect 63210 13530 63700 18150
rect 62740 13520 63700 13530
rect 49700 13380 63700 13520
rect 49690 13190 63700 13380
rect 49690 9010 49950 13190
rect 62740 13180 63700 13190
rect 53670 11120 53850 11130
rect 53850 10990 58640 11120
rect 53670 10980 53850 10990
rect 53680 10700 53820 10980
rect 49690 9000 49958 9010
rect 49690 8768 49958 8778
rect 49690 8760 49950 8768
rect 58480 4220 58640 10990
rect 92330 9590 92530 9600
rect 88510 9450 92330 9580
rect 64880 4320 67740 4430
rect 64450 4270 64620 4280
rect 26770 3980 27500 4130
rect 55560 4110 55750 4120
rect 53610 3940 55560 4110
rect 53610 3630 53780 3940
rect 55560 3930 55750 3940
rect 56220 4110 56410 4120
rect 56900 4110 57070 4120
rect 56410 3940 56900 4110
rect 57070 3940 58250 4110
rect 56220 3930 56410 3940
rect 56900 3930 57070 3940
rect 58080 3810 58250 3940
rect 58080 580 58250 3640
rect 58480 4050 64450 4220
rect 58480 950 58640 4050
rect 64450 4040 64620 4050
rect 64880 3810 65010 4320
rect 67590 4000 67740 4320
rect 67590 3830 67740 3840
rect 64880 3630 65010 3640
rect 78710 1810 78850 1820
rect 76930 1800 77050 1810
rect 75440 1600 75560 1610
rect 68130 1580 68240 1590
rect 68130 1400 68240 1410
rect 69920 1580 70040 1590
rect 69920 1400 70040 1410
rect 72110 1580 72360 1590
rect 72360 1410 73270 1580
rect 75440 1410 75560 1420
rect 76930 1580 77050 1700
rect 78710 1580 78850 1710
rect 76930 1430 77350 1580
rect 76930 1410 77100 1430
rect 78710 1410 79150 1580
rect 72110 1400 72360 1410
rect 58480 820 59010 950
rect 58080 430 58720 580
rect 43360 390 43600 400
rect 32030 -480 32270 -470
rect 32030 -10720 32270 -670
rect 41100 -1270 41300 -1260
rect 41100 -2860 41300 -1440
rect 41100 -3020 41300 -3010
rect 43360 -2860 43600 210
rect 45470 390 45760 400
rect 45470 200 45760 210
rect 43360 -3050 43600 -3040
rect 45490 -3150 45710 200
rect 58540 -1480 58720 430
rect 58190 -1630 58720 -1480
rect 45470 -3160 45740 -3150
rect 45470 -3380 45740 -3370
rect 58190 -8470 58350 -1630
rect 58850 -1880 59010 820
rect 88510 170 88650 9450
rect 92330 9440 92530 9450
rect 90520 9160 90790 9170
rect 90790 8930 92450 9160
rect 90520 8920 90790 8930
rect 80080 90 88650 170
rect 80080 80 88510 90
rect 75500 -800 75650 -790
rect 75500 -1040 75650 -1030
rect 58480 -2020 59010 -1880
rect 58480 -7220 58640 -2020
rect 73860 -2030 74050 -2020
rect 71770 -2040 71960 -2030
rect 71960 -2210 73860 -2040
rect 73860 -2220 74050 -2210
rect 71770 -2230 71960 -2220
rect 58480 -7350 59410 -7220
rect 58190 -8640 59090 -8470
rect 32030 -10880 59980 -10720
rect 32030 -10890 38240 -10880
<< via2 >>
rect 51800 18560 51980 18660
rect 52060 18560 52240 18660
rect 53670 10990 53850 11120
rect 55560 3940 55750 4110
rect 56220 3940 56410 4110
rect 56900 3940 57070 4110
rect 58080 3640 58250 3810
rect 64450 4050 64620 4270
rect 64880 3640 65010 3810
rect 76930 1700 77050 1800
rect 68130 1410 68240 1580
rect 69920 1410 70040 1580
rect 72110 1410 72360 1580
rect 75440 1420 75560 1600
rect 78710 1710 78850 1810
rect 43360 210 43600 390
rect 32030 -670 32270 -480
rect 41100 -1440 41300 -1270
rect 41100 -3010 41300 -2860
rect 45470 210 45760 390
rect 43360 -3040 43600 -2860
rect 45470 -3370 45740 -3160
rect 90520 8930 90790 9160
rect 75500 -1030 75650 -800
rect 71770 -2220 71960 -2040
rect 73860 -2210 74050 -2030
<< metal3 >>
rect 51790 18660 51990 18665
rect 51790 18560 51800 18660
rect 51980 18560 51990 18660
rect 51790 18555 51990 18560
rect 52050 18660 52250 18665
rect 52050 18560 52060 18660
rect 52240 18560 52250 18660
rect 52050 18555 52250 18560
rect 51840 14150 51970 18555
rect 52050 14400 52180 18555
rect 52050 14230 57070 14400
rect 51840 14020 53850 14150
rect 53670 11125 53850 14020
rect 53660 11120 53860 11125
rect 53660 10990 53670 11120
rect 53850 10990 53860 11120
rect 53660 10985 53860 10990
rect 25020 10260 28020 10360
rect 14700 -460 15020 -200
rect 25020 -460 25160 10260
rect 29000 10100 29140 10840
rect 26460 9980 29140 10100
rect 26460 600 26620 9980
rect 56900 4115 57070 14230
rect 90510 9160 90800 9165
rect 90510 8930 90520 9160
rect 90790 8930 90800 9160
rect 90510 8925 90800 8930
rect 64440 4270 65520 4330
rect 55550 4110 55760 4115
rect 56210 4110 56420 4115
rect 55550 3940 55560 4110
rect 55750 3940 56220 4110
rect 56410 3940 56420 4110
rect 55550 3935 55760 3940
rect 56210 3935 56420 3940
rect 56890 4110 57080 4115
rect 56890 3940 56900 4110
rect 57070 3940 57080 4110
rect 64440 4050 64450 4270
rect 64620 4220 65520 4270
rect 64620 4050 64630 4220
rect 65330 4080 65520 4220
rect 64440 4045 64630 4050
rect 56890 3935 57080 3940
rect 58070 3810 58260 3815
rect 64870 3810 65020 3815
rect 58070 3640 58080 3810
rect 58250 3640 64880 3810
rect 65010 3640 65020 3810
rect 58070 3635 58260 3640
rect 64870 3635 65020 3640
rect 29890 1080 30530 1240
rect 30360 660 30530 1080
rect 26460 460 27220 600
rect 30360 520 31690 660
rect 14700 -600 25160 -460
rect 31540 -1790 31690 520
rect 32030 -475 32270 1240
rect 33120 790 33470 1370
rect 33120 -160 33450 790
rect 34610 470 34840 1210
rect 34600 310 34610 470
rect 34840 310 34850 470
rect 36760 390 36990 1180
rect 36750 260 36760 390
rect 36990 260 37000 390
rect 38960 340 39190 1100
rect 41090 340 41320 1080
rect 43360 395 43590 1120
rect 45490 395 45720 1120
rect 43350 390 43610 395
rect 38950 210 38960 340
rect 39190 210 39200 340
rect 41080 210 41090 340
rect 41320 210 41330 340
rect 43350 210 43360 390
rect 43600 210 43610 390
rect 38960 180 39190 210
rect 41090 160 41320 210
rect 43350 205 43610 210
rect 45460 390 45770 395
rect 47710 390 47940 1120
rect 45460 210 45470 390
rect 45760 210 45770 390
rect 45460 205 45770 210
rect 43360 200 43590 205
rect 45490 200 45720 205
rect 47680 190 47690 390
rect 47950 190 47960 390
rect 33120 -380 33130 -160
rect 33450 -380 33460 -160
rect 33120 -410 33450 -380
rect 32020 -480 32280 -475
rect 32020 -670 32030 -480
rect 32270 -670 32280 -480
rect 32020 -675 32280 -670
rect 41090 -1270 41310 -1265
rect 41090 -1440 41100 -1270
rect 41300 -1440 41310 -1270
rect 41090 -1445 41310 -1440
rect 56630 -1790 57020 1940
rect 67470 1710 70050 1850
rect 78700 1810 78860 1815
rect 57940 390 57990 470
rect 31540 -2130 57020 -1790
rect 67470 -2300 67600 1710
rect 68120 1580 68250 1585
rect 32520 -2310 67600 -2300
rect 32520 -2440 36770 -2310
rect 36980 -2440 67600 -2310
rect 32520 -2460 67600 -2440
rect 67670 1410 68130 1580
rect 68240 1410 68250 1580
rect 67670 550 67820 1410
rect 68120 1405 68250 1410
rect 69910 1580 70050 1710
rect 76920 1800 77060 1805
rect 76920 1700 76930 1800
rect 77050 1700 77060 1800
rect 78700 1710 78710 1810
rect 78850 1710 78860 1810
rect 78700 1705 78860 1710
rect 76920 1695 77060 1700
rect 75430 1600 75570 1605
rect 69910 1410 69920 1580
rect 70040 1410 70050 1580
rect 69910 1405 70050 1410
rect 72100 1580 72370 1585
rect 72100 1410 72110 1580
rect 72360 1410 72370 1580
rect 75430 1420 75440 1600
rect 75560 1420 75570 1600
rect 75430 1415 75570 1420
rect 72100 1405 72370 1410
rect 67670 -2540 67800 550
rect 72760 -180 75380 -170
rect 72760 -310 76510 -180
rect 76650 -310 76660 -180
rect 72760 -320 75380 -310
rect 71760 -2040 71970 -2035
rect 71760 -2220 71770 -2040
rect 71960 -2220 71970 -2040
rect 71760 -2225 71970 -2220
rect 33370 -2550 67800 -2540
rect 33370 -2690 34620 -2550
rect 34830 -2690 67800 -2550
rect 33370 -2700 67800 -2690
rect 72760 -2850 72950 -320
rect 41090 -2860 41310 -2855
rect 41090 -3010 41100 -2860
rect 41300 -3010 41310 -2860
rect 43350 -2860 43610 -2855
rect 43350 -2880 43360 -2860
rect 41090 -3015 41310 -3010
rect 41580 -3040 43360 -2880
rect 43600 -2880 43610 -2860
rect 56520 -2870 72950 -2850
rect 56490 -2880 72950 -2870
rect 43600 -3040 72950 -2880
rect 73030 -570 78380 -440
rect 78530 -570 78540 -440
rect 43350 -3045 43610 -3040
rect 45460 -3160 45750 -3155
rect 73030 -3160 73190 -570
rect 75450 -795 75650 -790
rect 75450 -800 75660 -795
rect 75450 -1030 75500 -800
rect 75650 -1030 75660 -800
rect 75450 -1035 75660 -1030
rect 73850 -2030 74060 -2025
rect 73850 -2210 73860 -2030
rect 74050 -2210 74060 -2030
rect 73850 -2215 74060 -2210
rect 75450 -3160 75650 -1035
rect 45460 -3180 45470 -3160
rect 41580 -3340 45470 -3180
rect 44790 -3350 45470 -3340
rect 45460 -3370 45470 -3350
rect 45740 -3180 45750 -3160
rect 45740 -3190 47420 -3180
rect 56510 -3190 73190 -3160
rect 45740 -3350 73190 -3190
rect 75440 -3300 75450 -3160
rect 75650 -3300 75660 -3160
rect 45740 -3370 45750 -3350
rect 45460 -3375 45750 -3370
<< via3 >>
rect 90520 8930 90790 9160
rect 34610 310 34840 470
rect 36760 260 36990 390
rect 38960 210 39190 340
rect 41090 210 41320 340
rect 47690 190 47950 390
rect 33130 -380 33450 -160
rect 41100 -1440 41300 -1270
rect 36770 -2440 36980 -2310
rect 76930 1700 77050 1800
rect 78710 1710 78850 1810
rect 72110 1410 72360 1580
rect 75440 1420 75560 1600
rect 76510 -310 76650 -180
rect 71770 -2220 71960 -2040
rect 34620 -2690 34830 -2550
rect 41100 -3010 41300 -2860
rect 78380 -570 78530 -440
rect 73860 -2210 74050 -2030
rect 75450 -3300 75650 -3160
<< metal4 >>
rect 90519 9160 90791 9161
rect 90519 8930 90520 9160
rect 90790 8930 90791 9160
rect 90519 8929 90791 8930
rect 78709 1810 78851 1811
rect 76929 1800 77051 1801
rect 76929 1700 76930 1800
rect 77050 1700 77051 1800
rect 78709 1710 78710 1810
rect 78850 1710 78851 1810
rect 78709 1709 78851 1710
rect 76929 1699 77051 1700
rect 75439 1600 75561 1601
rect 72109 1580 72361 1581
rect 72109 1570 72110 1580
rect 72010 1410 72110 1570
rect 72360 1410 72361 1580
rect 75439 1570 75440 1600
rect 72010 1409 72361 1410
rect 73570 1420 75440 1570
rect 75560 1420 75561 1600
rect 76930 1560 77050 1699
rect 34609 470 34841 471
rect 34609 310 34610 470
rect 34840 310 34841 470
rect 34609 309 34841 310
rect 36759 390 36991 391
rect 33130 -159 33450 -130
rect 33129 -160 33451 -159
rect 33129 -380 33130 -160
rect 33450 -380 33451 -160
rect 33129 -381 33451 -380
rect 33130 -3120 33450 -381
rect 34610 -2550 34840 309
rect 36759 260 36760 390
rect 36990 260 36991 390
rect 38960 341 39190 410
rect 47689 390 47951 391
rect 41090 341 41320 380
rect 36759 259 36991 260
rect 38959 340 39191 341
rect 36760 -2310 36990 259
rect 38959 210 38960 340
rect 39190 210 39191 340
rect 38959 209 39191 210
rect 41089 340 41321 341
rect 41089 210 41090 340
rect 41320 210 41321 340
rect 41089 209 41321 210
rect 36760 -2440 36770 -2310
rect 36980 -2440 36990 -2310
rect 36760 -2460 36990 -2440
rect 34610 -2690 34620 -2550
rect 34830 -2690 34840 -2550
rect 34610 -2700 34840 -2690
rect 38960 -2590 39190 209
rect 41090 -1270 41320 209
rect 47689 190 47690 390
rect 47950 330 47951 390
rect 47950 190 47960 330
rect 47689 189 47960 190
rect 41090 -1440 41100 -1270
rect 41300 -1440 41320 -1270
rect 41090 -1460 41320 -1440
rect 47700 -2040 47960 189
rect 62480 -60 64200 -10
rect 62480 -890 63630 -60
rect 72010 -220 72170 1409
rect 72010 -340 72490 -220
rect 62480 -930 64200 -890
rect 71769 -2040 71961 -2039
rect 47700 -2220 71770 -2040
rect 71960 -2220 71961 -2040
rect 47700 -2230 47960 -2220
rect 71769 -2221 71961 -2220
rect 38960 -2600 56810 -2590
rect 72280 -2600 72490 -340
rect 38960 -2750 72490 -2600
rect 38960 -2760 56810 -2750
rect 41090 -2860 59740 -2850
rect 41090 -3010 41100 -2860
rect 41300 -2870 59740 -2860
rect 73570 -2870 73710 1420
rect 75439 1419 75561 1420
rect 76510 1450 77050 1560
rect 78710 1490 78850 1709
rect 76510 -179 76650 1450
rect 76930 1400 77050 1450
rect 78380 1380 78850 1490
rect 76509 -180 76651 -179
rect 76509 -310 76510 -180
rect 76650 -310 76651 -180
rect 76509 -311 76651 -310
rect 78380 -439 78530 1380
rect 78379 -440 78531 -439
rect 78379 -570 78380 -440
rect 78530 -570 78531 -440
rect 78379 -571 78531 -570
rect 90520 -2000 90790 8929
rect 73859 -2030 74051 -2029
rect 75930 -2030 90830 -2000
rect 73859 -2210 73860 -2030
rect 74050 -2200 90830 -2030
rect 74050 -2210 74051 -2200
rect 73859 -2211 74051 -2210
rect 41300 -3010 73710 -2870
rect 41090 -3020 73710 -3010
rect 33120 -3130 45770 -3120
rect 33120 -3150 59430 -3130
rect 33120 -3160 75700 -3150
rect 33120 -3300 75450 -3160
rect 75650 -3300 75700 -3160
rect 75449 -3301 75651 -3300
<< via4 >>
rect 63630 -890 64270 -60
<< metal5 >>
rect -1500 29120 136780 32790
rect 37900 12540 40060 29120
rect 50860 23600 52120 29120
rect 36860 12180 40060 12540
rect 25380 9300 28020 9760
rect 37900 9440 40060 12180
rect 49030 13540 49770 14890
rect 49030 10250 49760 13540
rect 15420 -1700 16220 -260
rect 16620 -600 17420 -180
rect 25380 -600 26100 9300
rect 49240 8750 49760 10250
rect 66360 9040 67460 29120
rect 16620 -1320 26100 -600
rect 27040 -1700 28640 -1020
rect 15420 -2320 28640 -1700
rect 45780 -2000 47800 -1020
rect 49030 -2000 49760 8750
rect 62400 7620 67460 9040
rect 66360 4220 67460 7620
rect 63640 -36 64290 10
rect 63606 -60 64294 -36
rect 63606 -890 63630 -60
rect 64270 -890 64294 -60
rect 63606 -914 64294 -890
rect 55510 -2000 59210 -1990
rect 61236 -2000 62204 -1976
rect 63640 -2000 64290 -914
rect 74560 -2000 75080 -960
rect 45780 -2350 75120 -2000
rect 45780 -20350 47800 -2350
rect 61236 -2404 62204 -2350
rect 83280 -3840 88000 29120
rect 112580 -1090 141180 440
rect 83020 -20350 88220 -18340
rect -1470 -21060 136810 -20350
rect 139420 -21060 141100 -1090
rect -1470 -22860 141290 -21060
rect -1470 -24020 136810 -22860
use comparator  comparator_0 ~/code/particle_detector/mag/comp
timestamp 1654768133
transform 1 0 74820 0 1 964
box -9660 -2484 5770 3520
use curr_mirror_channel  curr_mirror_channel_0 ~/code/particle_detector/mag/bias
timestamp 1654768133
transform 1 0 27070 0 1 -1680
box -20 0 21830 11434
use curr_mirror_distribution  curr_mirror_distribution_0 ~/code/particle_detector/mag/bias
timestamp 1654768133
transform 1 0 27190 0 1 10240
box 0 0 9830 2300
use fb_dark_current  fb_dark_current_0 ~/code/particle_detector/mag/feedback
timestamp 1654768133
transform 1 0 50550 0 1 16570
box -7920 -2510 12812 7750
use isource  isource_0 ~/code/particle_detector/mag/isource
timestamp 1654768133
transform 1 0 -180 0 1 4490
box -280 -4830 23120 15920
use outd  outd_0 ~/code/particle_detector/mag/outd
timestamp 1654768133
transform 1 0 80030 0 1 -18650
box -30220 -60 57040 15224
use tia_core  tia_core_0 ~/code/particle_detector/mag/tia
timestamp 1654768133
transform 1 0 51540 0 1 10030
box -1860 -11680 11730 2790
use transmitter  transmitter_0 ~/code/particle_detector/mag/lvds
timestamp 1654771420
transform 1 0 92230 0 1 5554
box -10 -6994 21080 20114
<< labels >>
rlabel metal5 -610 -23380 1100 -21480 1 VN
rlabel metal5 -30 30358 1770 31878 1 VP_an
rlabel metal2 49800 13250 50120 13480 1 In_Tia
rlabel metal3 57940 390 57990 470 1 Dis_TIA
rlabel metal1 49550 14950 49610 14980 1 Dis_Feedback
rlabel metal3 33150 50 33370 200 1 ctl_bias
rlabel metal4 34650 90 34790 270 1 comp_bias_1
rlabel metal4 36810 70 36950 250 1 comp_bias_2
rlabel metal4 38990 -10 39130 170 1 comp_bias_3
rlabel metal4 41110 -60 41250 120 1 comp_bias_4
rlabel metal2 45520 20 45650 140 1 comp_bias_6
rlabel metal2 43390 -20 43550 130 1 comp_bias_5
rlabel metal4 47740 -130 47900 20 1 bias_lvds
<< end >>
