magic
tech sky130A
magscale 1 2
timestamp 1645787783
<< error_p >>
rect -1107 272 -1049 278
rect -911 272 -853 278
rect -715 272 -657 278
rect -519 272 -461 278
rect -323 272 -265 278
rect -127 272 -69 278
rect 69 272 127 278
rect 265 272 323 278
rect 461 272 519 278
rect 657 272 715 278
rect 853 272 911 278
rect 1049 272 1107 278
rect -1107 238 -1095 272
rect -911 238 -899 272
rect -715 238 -703 272
rect -519 238 -507 272
rect -323 238 -311 272
rect -127 238 -115 272
rect 69 238 81 272
rect 265 238 277 272
rect 461 238 473 272
rect 657 238 669 272
rect 853 238 865 272
rect 1049 238 1061 272
rect -1107 232 -1049 238
rect -911 232 -853 238
rect -715 232 -657 238
rect -519 232 -461 238
rect -323 232 -265 238
rect -127 232 -69 238
rect 69 232 127 238
rect 265 232 323 238
rect 461 232 519 238
rect 657 232 715 238
rect 853 232 911 238
rect 1049 232 1107 238
rect -1205 -238 -1147 -232
rect -1009 -238 -951 -232
rect -813 -238 -755 -232
rect -617 -238 -559 -232
rect -421 -238 -363 -232
rect -225 -238 -167 -232
rect -29 -238 29 -232
rect 167 -238 225 -232
rect 363 -238 421 -232
rect 559 -238 617 -232
rect 755 -238 813 -232
rect 951 -238 1009 -232
rect 1147 -238 1205 -232
rect -1205 -272 -1193 -238
rect -1009 -272 -997 -238
rect -813 -272 -801 -238
rect -617 -272 -605 -238
rect -421 -272 -409 -238
rect -225 -272 -213 -238
rect -29 -272 -17 -238
rect 167 -272 179 -238
rect 363 -272 375 -238
rect 559 -272 571 -238
rect 755 -272 767 -238
rect 951 -272 963 -238
rect 1147 -272 1159 -238
rect -1205 -278 -1147 -272
rect -1009 -278 -951 -272
rect -813 -278 -755 -272
rect -617 -278 -559 -272
rect -421 -278 -363 -272
rect -225 -278 -167 -272
rect -29 -278 29 -272
rect 167 -278 225 -272
rect 363 -278 421 -272
rect 559 -278 617 -272
rect 755 -278 813 -272
rect 951 -278 1009 -272
rect 1147 -278 1205 -272
<< pwell >>
rect -1392 -410 1392 410
<< nmos >>
rect -1196 -200 -1156 200
rect -1098 -200 -1058 200
rect -1000 -200 -960 200
rect -902 -200 -862 200
rect -804 -200 -764 200
rect -706 -200 -666 200
rect -608 -200 -568 200
rect -510 -200 -470 200
rect -412 -200 -372 200
rect -314 -200 -274 200
rect -216 -200 -176 200
rect -118 -200 -78 200
rect -20 -200 20 200
rect 78 -200 118 200
rect 176 -200 216 200
rect 274 -200 314 200
rect 372 -200 412 200
rect 470 -200 510 200
rect 568 -200 608 200
rect 666 -200 706 200
rect 764 -200 804 200
rect 862 -200 902 200
rect 960 -200 1000 200
rect 1058 -200 1098 200
rect 1156 -200 1196 200
<< ndiff >>
rect -1254 188 -1196 200
rect -1254 -188 -1242 188
rect -1208 -188 -1196 188
rect -1254 -200 -1196 -188
rect -1156 188 -1098 200
rect -1156 -188 -1144 188
rect -1110 -188 -1098 188
rect -1156 -200 -1098 -188
rect -1058 188 -1000 200
rect -1058 -188 -1046 188
rect -1012 -188 -1000 188
rect -1058 -200 -1000 -188
rect -960 188 -902 200
rect -960 -188 -948 188
rect -914 -188 -902 188
rect -960 -200 -902 -188
rect -862 188 -804 200
rect -862 -188 -850 188
rect -816 -188 -804 188
rect -862 -200 -804 -188
rect -764 188 -706 200
rect -764 -188 -752 188
rect -718 -188 -706 188
rect -764 -200 -706 -188
rect -666 188 -608 200
rect -666 -188 -654 188
rect -620 -188 -608 188
rect -666 -200 -608 -188
rect -568 188 -510 200
rect -568 -188 -556 188
rect -522 -188 -510 188
rect -568 -200 -510 -188
rect -470 188 -412 200
rect -470 -188 -458 188
rect -424 -188 -412 188
rect -470 -200 -412 -188
rect -372 188 -314 200
rect -372 -188 -360 188
rect -326 -188 -314 188
rect -372 -200 -314 -188
rect -274 188 -216 200
rect -274 -188 -262 188
rect -228 -188 -216 188
rect -274 -200 -216 -188
rect -176 188 -118 200
rect -176 -188 -164 188
rect -130 -188 -118 188
rect -176 -200 -118 -188
rect -78 188 -20 200
rect -78 -188 -66 188
rect -32 -188 -20 188
rect -78 -200 -20 -188
rect 20 188 78 200
rect 20 -188 32 188
rect 66 -188 78 188
rect 20 -200 78 -188
rect 118 188 176 200
rect 118 -188 130 188
rect 164 -188 176 188
rect 118 -200 176 -188
rect 216 188 274 200
rect 216 -188 228 188
rect 262 -188 274 188
rect 216 -200 274 -188
rect 314 188 372 200
rect 314 -188 326 188
rect 360 -188 372 188
rect 314 -200 372 -188
rect 412 188 470 200
rect 412 -188 424 188
rect 458 -188 470 188
rect 412 -200 470 -188
rect 510 188 568 200
rect 510 -188 522 188
rect 556 -188 568 188
rect 510 -200 568 -188
rect 608 188 666 200
rect 608 -188 620 188
rect 654 -188 666 188
rect 608 -200 666 -188
rect 706 188 764 200
rect 706 -188 718 188
rect 752 -188 764 188
rect 706 -200 764 -188
rect 804 188 862 200
rect 804 -188 816 188
rect 850 -188 862 188
rect 804 -200 862 -188
rect 902 188 960 200
rect 902 -188 914 188
rect 948 -188 960 188
rect 902 -200 960 -188
rect 1000 188 1058 200
rect 1000 -188 1012 188
rect 1046 -188 1058 188
rect 1000 -200 1058 -188
rect 1098 188 1156 200
rect 1098 -188 1110 188
rect 1144 -188 1156 188
rect 1098 -200 1156 -188
rect 1196 188 1254 200
rect 1196 -188 1208 188
rect 1242 -188 1254 188
rect 1196 -200 1254 -188
<< ndiffc >>
rect -1242 -188 -1208 188
rect -1144 -188 -1110 188
rect -1046 -188 -1012 188
rect -948 -188 -914 188
rect -850 -188 -816 188
rect -752 -188 -718 188
rect -654 -188 -620 188
rect -556 -188 -522 188
rect -458 -188 -424 188
rect -360 -188 -326 188
rect -262 -188 -228 188
rect -164 -188 -130 188
rect -66 -188 -32 188
rect 32 -188 66 188
rect 130 -188 164 188
rect 228 -188 262 188
rect 326 -188 360 188
rect 424 -188 458 188
rect 522 -188 556 188
rect 620 -188 654 188
rect 718 -188 752 188
rect 816 -188 850 188
rect 914 -188 948 188
rect 1012 -188 1046 188
rect 1110 -188 1144 188
rect 1208 -188 1242 188
<< psubdiff >>
rect -1356 340 -1260 374
rect 1260 340 1356 374
rect -1356 278 -1322 340
rect 1322 278 1356 340
rect -1356 -340 -1322 -278
rect 1322 -340 1356 -278
rect -1356 -374 -1260 -340
rect 1260 -374 1356 -340
<< psubdiffcont >>
rect -1260 340 1260 374
rect -1356 -278 -1322 278
rect 1322 -278 1356 278
rect -1260 -374 1260 -340
<< poly >>
rect -1111 272 -1045 288
rect -1111 238 -1095 272
rect -1061 238 -1045 272
rect -1196 200 -1156 226
rect -1111 222 -1045 238
rect -915 272 -849 288
rect -915 238 -899 272
rect -865 238 -849 272
rect -1098 200 -1058 222
rect -1000 200 -960 226
rect -915 222 -849 238
rect -719 272 -653 288
rect -719 238 -703 272
rect -669 238 -653 272
rect -902 200 -862 222
rect -804 200 -764 226
rect -719 222 -653 238
rect -523 272 -457 288
rect -523 238 -507 272
rect -473 238 -457 272
rect -706 200 -666 222
rect -608 200 -568 226
rect -523 222 -457 238
rect -327 272 -261 288
rect -327 238 -311 272
rect -277 238 -261 272
rect -510 200 -470 222
rect -412 200 -372 226
rect -327 222 -261 238
rect -131 272 -65 288
rect -131 238 -115 272
rect -81 238 -65 272
rect -314 200 -274 222
rect -216 200 -176 226
rect -131 222 -65 238
rect 65 272 131 288
rect 65 238 81 272
rect 115 238 131 272
rect -118 200 -78 222
rect -20 200 20 226
rect 65 222 131 238
rect 261 272 327 288
rect 261 238 277 272
rect 311 238 327 272
rect 78 200 118 222
rect 176 200 216 226
rect 261 222 327 238
rect 457 272 523 288
rect 457 238 473 272
rect 507 238 523 272
rect 274 200 314 222
rect 372 200 412 226
rect 457 222 523 238
rect 653 272 719 288
rect 653 238 669 272
rect 703 238 719 272
rect 470 200 510 222
rect 568 200 608 226
rect 653 222 719 238
rect 849 272 915 288
rect 849 238 865 272
rect 899 238 915 272
rect 666 200 706 222
rect 764 200 804 226
rect 849 222 915 238
rect 1045 272 1111 288
rect 1045 238 1061 272
rect 1095 238 1111 272
rect 862 200 902 222
rect 960 200 1000 226
rect 1045 222 1111 238
rect 1058 200 1098 222
rect 1156 200 1196 226
rect -1196 -222 -1156 -200
rect -1209 -238 -1143 -222
rect -1098 -226 -1058 -200
rect -1000 -222 -960 -200
rect -1209 -272 -1193 -238
rect -1159 -272 -1143 -238
rect -1209 -288 -1143 -272
rect -1013 -238 -947 -222
rect -902 -226 -862 -200
rect -804 -222 -764 -200
rect -1013 -272 -997 -238
rect -963 -272 -947 -238
rect -1013 -288 -947 -272
rect -817 -238 -751 -222
rect -706 -226 -666 -200
rect -608 -222 -568 -200
rect -817 -272 -801 -238
rect -767 -272 -751 -238
rect -817 -288 -751 -272
rect -621 -238 -555 -222
rect -510 -226 -470 -200
rect -412 -222 -372 -200
rect -621 -272 -605 -238
rect -571 -272 -555 -238
rect -621 -288 -555 -272
rect -425 -238 -359 -222
rect -314 -226 -274 -200
rect -216 -222 -176 -200
rect -425 -272 -409 -238
rect -375 -272 -359 -238
rect -425 -288 -359 -272
rect -229 -238 -163 -222
rect -118 -226 -78 -200
rect -20 -222 20 -200
rect -229 -272 -213 -238
rect -179 -272 -163 -238
rect -229 -288 -163 -272
rect -33 -238 33 -222
rect 78 -226 118 -200
rect 176 -222 216 -200
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
rect 163 -238 229 -222
rect 274 -226 314 -200
rect 372 -222 412 -200
rect 163 -272 179 -238
rect 213 -272 229 -238
rect 163 -288 229 -272
rect 359 -238 425 -222
rect 470 -226 510 -200
rect 568 -222 608 -200
rect 359 -272 375 -238
rect 409 -272 425 -238
rect 359 -288 425 -272
rect 555 -238 621 -222
rect 666 -226 706 -200
rect 764 -222 804 -200
rect 555 -272 571 -238
rect 605 -272 621 -238
rect 555 -288 621 -272
rect 751 -238 817 -222
rect 862 -226 902 -200
rect 960 -222 1000 -200
rect 751 -272 767 -238
rect 801 -272 817 -238
rect 751 -288 817 -272
rect 947 -238 1013 -222
rect 1058 -226 1098 -200
rect 1156 -222 1196 -200
rect 947 -272 963 -238
rect 997 -272 1013 -238
rect 947 -288 1013 -272
rect 1143 -238 1209 -222
rect 1143 -272 1159 -238
rect 1193 -272 1209 -238
rect 1143 -288 1209 -272
<< polycont >>
rect -1095 238 -1061 272
rect -899 238 -865 272
rect -703 238 -669 272
rect -507 238 -473 272
rect -311 238 -277 272
rect -115 238 -81 272
rect 81 238 115 272
rect 277 238 311 272
rect 473 238 507 272
rect 669 238 703 272
rect 865 238 899 272
rect 1061 238 1095 272
rect -1193 -272 -1159 -238
rect -997 -272 -963 -238
rect -801 -272 -767 -238
rect -605 -272 -571 -238
rect -409 -272 -375 -238
rect -213 -272 -179 -238
rect -17 -272 17 -238
rect 179 -272 213 -238
rect 375 -272 409 -238
rect 571 -272 605 -238
rect 767 -272 801 -238
rect 963 -272 997 -238
rect 1159 -272 1193 -238
<< locali >>
rect -1356 340 -1260 374
rect 1260 340 1356 374
rect -1356 278 -1322 340
rect 1322 278 1356 340
rect -1111 238 -1095 272
rect -1061 238 -1045 272
rect -915 238 -899 272
rect -865 238 -849 272
rect -719 238 -703 272
rect -669 238 -653 272
rect -523 238 -507 272
rect -473 238 -457 272
rect -327 238 -311 272
rect -277 238 -261 272
rect -131 238 -115 272
rect -81 238 -65 272
rect 65 238 81 272
rect 115 238 131 272
rect 261 238 277 272
rect 311 238 327 272
rect 457 238 473 272
rect 507 238 523 272
rect 653 238 669 272
rect 703 238 719 272
rect 849 238 865 272
rect 899 238 915 272
rect 1045 238 1061 272
rect 1095 238 1111 272
rect -1242 188 -1208 204
rect -1242 -204 -1208 -188
rect -1144 188 -1110 204
rect -1144 -204 -1110 -188
rect -1046 188 -1012 204
rect -1046 -204 -1012 -188
rect -948 188 -914 204
rect -948 -204 -914 -188
rect -850 188 -816 204
rect -850 -204 -816 -188
rect -752 188 -718 204
rect -752 -204 -718 -188
rect -654 188 -620 204
rect -654 -204 -620 -188
rect -556 188 -522 204
rect -556 -204 -522 -188
rect -458 188 -424 204
rect -458 -204 -424 -188
rect -360 188 -326 204
rect -360 -204 -326 -188
rect -262 188 -228 204
rect -262 -204 -228 -188
rect -164 188 -130 204
rect -164 -204 -130 -188
rect -66 188 -32 204
rect -66 -204 -32 -188
rect 32 188 66 204
rect 32 -204 66 -188
rect 130 188 164 204
rect 130 -204 164 -188
rect 228 188 262 204
rect 228 -204 262 -188
rect 326 188 360 204
rect 326 -204 360 -188
rect 424 188 458 204
rect 424 -204 458 -188
rect 522 188 556 204
rect 522 -204 556 -188
rect 620 188 654 204
rect 620 -204 654 -188
rect 718 188 752 204
rect 718 -204 752 -188
rect 816 188 850 204
rect 816 -204 850 -188
rect 914 188 948 204
rect 914 -204 948 -188
rect 1012 188 1046 204
rect 1012 -204 1046 -188
rect 1110 188 1144 204
rect 1110 -204 1144 -188
rect 1208 188 1242 204
rect 1208 -204 1242 -188
rect -1209 -272 -1193 -238
rect -1159 -272 -1143 -238
rect -1013 -272 -997 -238
rect -963 -272 -947 -238
rect -817 -272 -801 -238
rect -767 -272 -751 -238
rect -621 -272 -605 -238
rect -571 -272 -555 -238
rect -425 -272 -409 -238
rect -375 -272 -359 -238
rect -229 -272 -213 -238
rect -179 -272 -163 -238
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 163 -272 179 -238
rect 213 -272 229 -238
rect 359 -272 375 -238
rect 409 -272 425 -238
rect 555 -272 571 -238
rect 605 -272 621 -238
rect 751 -272 767 -238
rect 801 -272 817 -238
rect 947 -272 963 -238
rect 997 -272 1013 -238
rect 1143 -272 1159 -238
rect 1193 -272 1209 -238
rect -1356 -340 -1322 -278
rect 1322 -340 1356 -278
rect -1356 -374 -1260 -340
rect 1260 -374 1356 -340
<< viali >>
rect -1095 238 -1061 272
rect -899 238 -865 272
rect -703 238 -669 272
rect -507 238 -473 272
rect -311 238 -277 272
rect -115 238 -81 272
rect 81 238 115 272
rect 277 238 311 272
rect 473 238 507 272
rect 669 238 703 272
rect 865 238 899 272
rect 1061 238 1095 272
rect -1242 -188 -1208 188
rect -1144 -188 -1110 188
rect -1046 -188 -1012 188
rect -948 -188 -914 188
rect -850 -188 -816 188
rect -752 -188 -718 188
rect -654 -188 -620 188
rect -556 -188 -522 188
rect -458 -188 -424 188
rect -360 -188 -326 188
rect -262 -188 -228 188
rect -164 -188 -130 188
rect -66 -188 -32 188
rect 32 -188 66 188
rect 130 -188 164 188
rect 228 -188 262 188
rect 326 -188 360 188
rect 424 -188 458 188
rect 522 -188 556 188
rect 620 -188 654 188
rect 718 -188 752 188
rect 816 -188 850 188
rect 914 -188 948 188
rect 1012 -188 1046 188
rect 1110 -188 1144 188
rect 1208 -188 1242 188
rect -1193 -272 -1159 -238
rect -997 -272 -963 -238
rect -801 -272 -767 -238
rect -605 -272 -571 -238
rect -409 -272 -375 -238
rect -213 -272 -179 -238
rect -17 -272 17 -238
rect 179 -272 213 -238
rect 375 -272 409 -238
rect 571 -272 605 -238
rect 767 -272 801 -238
rect 963 -272 997 -238
rect 1159 -272 1193 -238
<< metal1 >>
rect -1107 272 -1049 278
rect -1107 238 -1095 272
rect -1061 238 -1049 272
rect -1107 232 -1049 238
rect -911 272 -853 278
rect -911 238 -899 272
rect -865 238 -853 272
rect -911 232 -853 238
rect -715 272 -657 278
rect -715 238 -703 272
rect -669 238 -657 272
rect -715 232 -657 238
rect -519 272 -461 278
rect -519 238 -507 272
rect -473 238 -461 272
rect -519 232 -461 238
rect -323 272 -265 278
rect -323 238 -311 272
rect -277 238 -265 272
rect -323 232 -265 238
rect -127 272 -69 278
rect -127 238 -115 272
rect -81 238 -69 272
rect -127 232 -69 238
rect 69 272 127 278
rect 69 238 81 272
rect 115 238 127 272
rect 69 232 127 238
rect 265 272 323 278
rect 265 238 277 272
rect 311 238 323 272
rect 265 232 323 238
rect 461 272 519 278
rect 461 238 473 272
rect 507 238 519 272
rect 461 232 519 238
rect 657 272 715 278
rect 657 238 669 272
rect 703 238 715 272
rect 657 232 715 238
rect 853 272 911 278
rect 853 238 865 272
rect 899 238 911 272
rect 853 232 911 238
rect 1049 272 1107 278
rect 1049 238 1061 272
rect 1095 238 1107 272
rect 1049 232 1107 238
rect -1248 188 -1202 200
rect -1248 -188 -1242 188
rect -1208 -188 -1202 188
rect -1248 -200 -1202 -188
rect -1150 188 -1104 200
rect -1150 -188 -1144 188
rect -1110 -188 -1104 188
rect -1150 -200 -1104 -188
rect -1052 188 -1006 200
rect -1052 -188 -1046 188
rect -1012 -188 -1006 188
rect -1052 -200 -1006 -188
rect -954 188 -908 200
rect -954 -188 -948 188
rect -914 -188 -908 188
rect -954 -200 -908 -188
rect -856 188 -810 200
rect -856 -188 -850 188
rect -816 -188 -810 188
rect -856 -200 -810 -188
rect -758 188 -712 200
rect -758 -188 -752 188
rect -718 -188 -712 188
rect -758 -200 -712 -188
rect -660 188 -614 200
rect -660 -188 -654 188
rect -620 -188 -614 188
rect -660 -200 -614 -188
rect -562 188 -516 200
rect -562 -188 -556 188
rect -522 -188 -516 188
rect -562 -200 -516 -188
rect -464 188 -418 200
rect -464 -188 -458 188
rect -424 -188 -418 188
rect -464 -200 -418 -188
rect -366 188 -320 200
rect -366 -188 -360 188
rect -326 -188 -320 188
rect -366 -200 -320 -188
rect -268 188 -222 200
rect -268 -188 -262 188
rect -228 -188 -222 188
rect -268 -200 -222 -188
rect -170 188 -124 200
rect -170 -188 -164 188
rect -130 -188 -124 188
rect -170 -200 -124 -188
rect -72 188 -26 200
rect -72 -188 -66 188
rect -32 -188 -26 188
rect -72 -200 -26 -188
rect 26 188 72 200
rect 26 -188 32 188
rect 66 -188 72 188
rect 26 -200 72 -188
rect 124 188 170 200
rect 124 -188 130 188
rect 164 -188 170 188
rect 124 -200 170 -188
rect 222 188 268 200
rect 222 -188 228 188
rect 262 -188 268 188
rect 222 -200 268 -188
rect 320 188 366 200
rect 320 -188 326 188
rect 360 -188 366 188
rect 320 -200 366 -188
rect 418 188 464 200
rect 418 -188 424 188
rect 458 -188 464 188
rect 418 -200 464 -188
rect 516 188 562 200
rect 516 -188 522 188
rect 556 -188 562 188
rect 516 -200 562 -188
rect 614 188 660 200
rect 614 -188 620 188
rect 654 -188 660 188
rect 614 -200 660 -188
rect 712 188 758 200
rect 712 -188 718 188
rect 752 -188 758 188
rect 712 -200 758 -188
rect 810 188 856 200
rect 810 -188 816 188
rect 850 -188 856 188
rect 810 -200 856 -188
rect 908 188 954 200
rect 908 -188 914 188
rect 948 -188 954 188
rect 908 -200 954 -188
rect 1006 188 1052 200
rect 1006 -188 1012 188
rect 1046 -188 1052 188
rect 1006 -200 1052 -188
rect 1104 188 1150 200
rect 1104 -188 1110 188
rect 1144 -188 1150 188
rect 1104 -200 1150 -188
rect 1202 188 1248 200
rect 1202 -188 1208 188
rect 1242 -188 1248 188
rect 1202 -200 1248 -188
rect -1205 -238 -1147 -232
rect -1205 -272 -1193 -238
rect -1159 -272 -1147 -238
rect -1205 -278 -1147 -272
rect -1009 -238 -951 -232
rect -1009 -272 -997 -238
rect -963 -272 -951 -238
rect -1009 -278 -951 -272
rect -813 -238 -755 -232
rect -813 -272 -801 -238
rect -767 -272 -755 -238
rect -813 -278 -755 -272
rect -617 -238 -559 -232
rect -617 -272 -605 -238
rect -571 -272 -559 -238
rect -617 -278 -559 -272
rect -421 -238 -363 -232
rect -421 -272 -409 -238
rect -375 -272 -363 -238
rect -421 -278 -363 -272
rect -225 -238 -167 -232
rect -225 -272 -213 -238
rect -179 -272 -167 -238
rect -225 -278 -167 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 167 -238 225 -232
rect 167 -272 179 -238
rect 213 -272 225 -238
rect 167 -278 225 -272
rect 363 -238 421 -232
rect 363 -272 375 -238
rect 409 -272 421 -238
rect 363 -278 421 -272
rect 559 -238 617 -232
rect 559 -272 571 -238
rect 605 -272 617 -238
rect 559 -278 617 -272
rect 755 -238 813 -232
rect 755 -272 767 -238
rect 801 -272 813 -238
rect 755 -278 813 -272
rect 951 -238 1009 -232
rect 951 -272 963 -238
rect 997 -272 1009 -238
rect 951 -278 1009 -272
rect 1147 -238 1205 -232
rect 1147 -272 1159 -238
rect 1193 -272 1205 -238
rect 1147 -278 1205 -272
<< properties >>
string FIXED_BBOX -1339 -357 1339 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.2 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
