magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< nwell >>
rect 132 600 870 666
rect 150 590 180 600
rect 342 590 372 600
rect 534 590 564 600
rect 726 592 756 600
rect 246 138 276 152
rect 438 138 468 152
rect 630 138 660 152
rect 822 138 852 152
rect 132 72 870 138
<< poly >>
rect 132 650 870 666
rect 132 616 148 650
rect 182 616 340 650
rect 374 616 532 650
rect 566 616 724 650
rect 758 616 870 650
rect 132 600 870 616
rect 150 590 180 600
rect 342 590 372 600
rect 534 590 564 600
rect 726 592 756 600
rect 246 138 276 152
rect 438 138 468 152
rect 630 138 660 152
rect 822 138 852 152
rect 132 122 870 138
rect 132 88 244 122
rect 278 88 436 122
rect 470 88 628 122
rect 662 88 820 122
rect 854 88 870 122
rect 132 72 870 88
<< polycont >>
rect 148 616 182 650
rect 340 616 374 650
rect 532 616 566 650
rect 724 616 758 650
rect 244 88 278 122
rect 436 88 470 122
rect 628 88 662 122
rect 820 88 854 122
<< locali >>
rect 10 830 110 1550
rect 440 830 540 1550
rect -10 740 560 820
rect 132 616 148 650
rect 182 616 340 650
rect 374 616 532 650
rect 566 616 724 650
rect 758 616 870 650
rect 132 88 244 122
rect 278 88 436 122
rect 470 88 628 122
rect 662 88 820 122
rect 854 88 870 122
<< viali >>
rect 148 616 182 650
rect 340 616 374 650
rect 532 616 566 650
rect 724 616 758 650
rect 244 88 278 122
rect 436 88 470 122
rect 628 88 662 122
rect 820 88 854 122
<< metal1 >>
rect 140 1430 580 1490
rect 70 1220 80 1390
rect 150 1220 160 1390
rect 390 1220 400 1390
rect 470 1220 480 1390
rect 230 990 240 1160
rect 310 990 320 1160
rect 520 950 580 1430
rect 140 890 580 950
rect 320 660 390 890
rect -10 650 870 660
rect -10 616 148 650
rect 182 616 340 650
rect 374 616 532 650
rect 566 616 724 650
rect 758 616 870 650
rect -10 610 870 616
rect -10 130 40 610
rect 80 400 90 570
rect 150 400 160 570
rect 270 400 280 570
rect 340 400 350 570
rect 460 400 470 570
rect 530 400 540 570
rect 650 400 660 570
rect 720 400 730 570
rect 850 400 860 570
rect 920 400 930 570
rect 170 170 180 340
rect 240 170 250 340
rect 370 170 380 340
rect 440 170 450 340
rect 560 170 570 340
rect 630 170 640 340
rect 750 170 760 340
rect 820 170 830 340
rect -10 122 870 130
rect -10 88 244 122
rect 278 88 436 122
rect 470 88 628 122
rect 662 88 820 122
rect 854 88 870 122
rect -10 80 870 88
<< via1 >>
rect 80 1220 150 1390
rect 400 1220 470 1390
rect 240 990 310 1160
rect 90 400 150 570
rect 280 400 340 570
rect 470 400 530 570
rect 660 400 720 570
rect 860 400 920 570
rect 180 170 240 340
rect 380 170 440 340
rect 570 170 630 340
rect 760 170 820 340
<< metal2 >>
rect 80 1390 150 1400
rect 400 1390 470 1400
rect 150 1220 400 1390
rect 80 1210 150 1220
rect 400 1210 470 1220
rect 240 1160 310 1170
rect 230 990 240 1160
rect 310 990 370 1160
rect 90 570 150 580
rect 230 570 370 990
rect 470 570 530 580
rect 660 570 720 580
rect 860 570 920 580
rect 150 400 280 570
rect 340 400 470 570
rect 530 400 660 570
rect 720 400 860 570
rect 90 390 150 400
rect 280 390 340 400
rect 470 390 530 400
rect 660 390 720 400
rect 860 390 920 400
rect 180 340 240 350
rect 380 340 440 350
rect 570 340 630 350
rect 760 340 820 350
rect 240 170 380 340
rect 440 170 570 340
rect 630 170 760 340
rect 180 160 240 170
rect 380 160 440 170
rect 570 160 630 170
rect 760 160 820 170
use sky130_fd_pr__pfet_01v8_PD4XN5  sky130_fd_pr__pfet_01v8_PD4XN5_0
timestamp 1654768133
transform 1 0 275 0 1 1189
box -325 -419 325 419
use sky130_fd_pr__pfet_01v8_U4PWGH  sky130_fd_pr__pfet_01v8_U4PWGH_0
timestamp 1654768133
transform 1 0 501 0 1 369
box -551 -419 551 419
<< end >>
