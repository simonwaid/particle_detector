magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< error_p >>
rect -557 1235 -499 1241
rect -365 1235 -307 1241
rect -173 1235 -115 1241
rect 19 1235 77 1241
rect 211 1235 269 1241
rect 403 1235 461 1241
rect -557 1201 -545 1235
rect -365 1201 -353 1235
rect -173 1201 -161 1235
rect 19 1201 31 1235
rect 211 1201 223 1235
rect 403 1201 415 1235
rect -557 1195 -499 1201
rect -365 1195 -307 1201
rect -173 1195 -115 1201
rect 19 1195 77 1201
rect 211 1195 269 1201
rect 403 1195 461 1201
rect -461 707 -403 713
rect -269 707 -211 713
rect -77 707 -19 713
rect 115 707 173 713
rect 307 707 365 713
rect 499 707 557 713
rect -461 673 -449 707
rect -269 673 -257 707
rect -77 673 -65 707
rect 115 673 127 707
rect 307 673 319 707
rect 499 673 511 707
rect -461 667 -403 673
rect -269 667 -211 673
rect -77 667 -19 673
rect 115 667 173 673
rect 307 667 365 673
rect 499 667 557 673
rect -461 599 -403 605
rect -269 599 -211 605
rect -77 599 -19 605
rect 115 599 173 605
rect 307 599 365 605
rect 499 599 557 605
rect -461 565 -449 599
rect -269 565 -257 599
rect -77 565 -65 599
rect 115 565 127 599
rect 307 565 319 599
rect 499 565 511 599
rect -461 559 -403 565
rect -269 559 -211 565
rect -77 559 -19 565
rect 115 559 173 565
rect 307 559 365 565
rect 499 559 557 565
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect -461 -565 -403 -559
rect -269 -565 -211 -559
rect -77 -565 -19 -559
rect 115 -565 173 -559
rect 307 -565 365 -559
rect 499 -565 557 -559
rect -461 -599 -449 -565
rect -269 -599 -257 -565
rect -77 -599 -65 -565
rect 115 -599 127 -565
rect 307 -599 319 -565
rect 499 -599 511 -565
rect -461 -605 -403 -599
rect -269 -605 -211 -599
rect -77 -605 -19 -599
rect 115 -605 173 -599
rect 307 -605 365 -599
rect 499 -605 557 -599
rect -461 -673 -403 -667
rect -269 -673 -211 -667
rect -77 -673 -19 -667
rect 115 -673 173 -667
rect 307 -673 365 -667
rect 499 -673 557 -667
rect -461 -707 -449 -673
rect -269 -707 -257 -673
rect -77 -707 -65 -673
rect 115 -707 127 -673
rect 307 -707 319 -673
rect 499 -707 511 -673
rect -461 -713 -403 -707
rect -269 -713 -211 -707
rect -77 -713 -19 -707
rect 115 -713 173 -707
rect 307 -713 365 -707
rect 499 -713 557 -707
rect -557 -1201 -499 -1195
rect -365 -1201 -307 -1195
rect -173 -1201 -115 -1195
rect 19 -1201 77 -1195
rect 211 -1201 269 -1195
rect 403 -1201 461 -1195
rect -557 -1235 -545 -1201
rect -365 -1235 -353 -1201
rect -173 -1235 -161 -1201
rect 19 -1235 31 -1201
rect 211 -1235 223 -1201
rect 403 -1235 415 -1201
rect -557 -1241 -499 -1235
rect -365 -1241 -307 -1235
rect -173 -1241 -115 -1235
rect 19 -1241 77 -1235
rect 211 -1241 269 -1235
rect 403 -1241 461 -1235
<< nwell >>
rect -743 -1373 743 1373
<< pmos >>
rect -543 754 -513 1154
rect -447 754 -417 1154
rect -351 754 -321 1154
rect -255 754 -225 1154
rect -159 754 -129 1154
rect -63 754 -33 1154
rect 33 754 63 1154
rect 129 754 159 1154
rect 225 754 255 1154
rect 321 754 351 1154
rect 417 754 447 1154
rect 513 754 543 1154
rect -543 118 -513 518
rect -447 118 -417 518
rect -351 118 -321 518
rect -255 118 -225 518
rect -159 118 -129 518
rect -63 118 -33 518
rect 33 118 63 518
rect 129 118 159 518
rect 225 118 255 518
rect 321 118 351 518
rect 417 118 447 518
rect 513 118 543 518
rect -543 -518 -513 -118
rect -447 -518 -417 -118
rect -351 -518 -321 -118
rect -255 -518 -225 -118
rect -159 -518 -129 -118
rect -63 -518 -33 -118
rect 33 -518 63 -118
rect 129 -518 159 -118
rect 225 -518 255 -118
rect 321 -518 351 -118
rect 417 -518 447 -118
rect 513 -518 543 -118
rect -543 -1154 -513 -754
rect -447 -1154 -417 -754
rect -351 -1154 -321 -754
rect -255 -1154 -225 -754
rect -159 -1154 -129 -754
rect -63 -1154 -33 -754
rect 33 -1154 63 -754
rect 129 -1154 159 -754
rect 225 -1154 255 -754
rect 321 -1154 351 -754
rect 417 -1154 447 -754
rect 513 -1154 543 -754
<< pdiff >>
rect -605 1142 -543 1154
rect -605 766 -593 1142
rect -559 766 -543 1142
rect -605 754 -543 766
rect -513 1142 -447 1154
rect -513 766 -497 1142
rect -463 766 -447 1142
rect -513 754 -447 766
rect -417 1142 -351 1154
rect -417 766 -401 1142
rect -367 766 -351 1142
rect -417 754 -351 766
rect -321 1142 -255 1154
rect -321 766 -305 1142
rect -271 766 -255 1142
rect -321 754 -255 766
rect -225 1142 -159 1154
rect -225 766 -209 1142
rect -175 766 -159 1142
rect -225 754 -159 766
rect -129 1142 -63 1154
rect -129 766 -113 1142
rect -79 766 -63 1142
rect -129 754 -63 766
rect -33 1142 33 1154
rect -33 766 -17 1142
rect 17 766 33 1142
rect -33 754 33 766
rect 63 1142 129 1154
rect 63 766 79 1142
rect 113 766 129 1142
rect 63 754 129 766
rect 159 1142 225 1154
rect 159 766 175 1142
rect 209 766 225 1142
rect 159 754 225 766
rect 255 1142 321 1154
rect 255 766 271 1142
rect 305 766 321 1142
rect 255 754 321 766
rect 351 1142 417 1154
rect 351 766 367 1142
rect 401 766 417 1142
rect 351 754 417 766
rect 447 1142 513 1154
rect 447 766 463 1142
rect 497 766 513 1142
rect 447 754 513 766
rect 543 1142 605 1154
rect 543 766 559 1142
rect 593 766 605 1142
rect 543 754 605 766
rect -605 506 -543 518
rect -605 130 -593 506
rect -559 130 -543 506
rect -605 118 -543 130
rect -513 506 -447 518
rect -513 130 -497 506
rect -463 130 -447 506
rect -513 118 -447 130
rect -417 506 -351 518
rect -417 130 -401 506
rect -367 130 -351 506
rect -417 118 -351 130
rect -321 506 -255 518
rect -321 130 -305 506
rect -271 130 -255 506
rect -321 118 -255 130
rect -225 506 -159 518
rect -225 130 -209 506
rect -175 130 -159 506
rect -225 118 -159 130
rect -129 506 -63 518
rect -129 130 -113 506
rect -79 130 -63 506
rect -129 118 -63 130
rect -33 506 33 518
rect -33 130 -17 506
rect 17 130 33 506
rect -33 118 33 130
rect 63 506 129 518
rect 63 130 79 506
rect 113 130 129 506
rect 63 118 129 130
rect 159 506 225 518
rect 159 130 175 506
rect 209 130 225 506
rect 159 118 225 130
rect 255 506 321 518
rect 255 130 271 506
rect 305 130 321 506
rect 255 118 321 130
rect 351 506 417 518
rect 351 130 367 506
rect 401 130 417 506
rect 351 118 417 130
rect 447 506 513 518
rect 447 130 463 506
rect 497 130 513 506
rect 447 118 513 130
rect 543 506 605 518
rect 543 130 559 506
rect 593 130 605 506
rect 543 118 605 130
rect -605 -130 -543 -118
rect -605 -506 -593 -130
rect -559 -506 -543 -130
rect -605 -518 -543 -506
rect -513 -130 -447 -118
rect -513 -506 -497 -130
rect -463 -506 -447 -130
rect -513 -518 -447 -506
rect -417 -130 -351 -118
rect -417 -506 -401 -130
rect -367 -506 -351 -130
rect -417 -518 -351 -506
rect -321 -130 -255 -118
rect -321 -506 -305 -130
rect -271 -506 -255 -130
rect -321 -518 -255 -506
rect -225 -130 -159 -118
rect -225 -506 -209 -130
rect -175 -506 -159 -130
rect -225 -518 -159 -506
rect -129 -130 -63 -118
rect -129 -506 -113 -130
rect -79 -506 -63 -130
rect -129 -518 -63 -506
rect -33 -130 33 -118
rect -33 -506 -17 -130
rect 17 -506 33 -130
rect -33 -518 33 -506
rect 63 -130 129 -118
rect 63 -506 79 -130
rect 113 -506 129 -130
rect 63 -518 129 -506
rect 159 -130 225 -118
rect 159 -506 175 -130
rect 209 -506 225 -130
rect 159 -518 225 -506
rect 255 -130 321 -118
rect 255 -506 271 -130
rect 305 -506 321 -130
rect 255 -518 321 -506
rect 351 -130 417 -118
rect 351 -506 367 -130
rect 401 -506 417 -130
rect 351 -518 417 -506
rect 447 -130 513 -118
rect 447 -506 463 -130
rect 497 -506 513 -130
rect 447 -518 513 -506
rect 543 -130 605 -118
rect 543 -506 559 -130
rect 593 -506 605 -130
rect 543 -518 605 -506
rect -605 -766 -543 -754
rect -605 -1142 -593 -766
rect -559 -1142 -543 -766
rect -605 -1154 -543 -1142
rect -513 -766 -447 -754
rect -513 -1142 -497 -766
rect -463 -1142 -447 -766
rect -513 -1154 -447 -1142
rect -417 -766 -351 -754
rect -417 -1142 -401 -766
rect -367 -1142 -351 -766
rect -417 -1154 -351 -1142
rect -321 -766 -255 -754
rect -321 -1142 -305 -766
rect -271 -1142 -255 -766
rect -321 -1154 -255 -1142
rect -225 -766 -159 -754
rect -225 -1142 -209 -766
rect -175 -1142 -159 -766
rect -225 -1154 -159 -1142
rect -129 -766 -63 -754
rect -129 -1142 -113 -766
rect -79 -1142 -63 -766
rect -129 -1154 -63 -1142
rect -33 -766 33 -754
rect -33 -1142 -17 -766
rect 17 -1142 33 -766
rect -33 -1154 33 -1142
rect 63 -766 129 -754
rect 63 -1142 79 -766
rect 113 -1142 129 -766
rect 63 -1154 129 -1142
rect 159 -766 225 -754
rect 159 -1142 175 -766
rect 209 -1142 225 -766
rect 159 -1154 225 -1142
rect 255 -766 321 -754
rect 255 -1142 271 -766
rect 305 -1142 321 -766
rect 255 -1154 321 -1142
rect 351 -766 417 -754
rect 351 -1142 367 -766
rect 401 -1142 417 -766
rect 351 -1154 417 -1142
rect 447 -766 513 -754
rect 447 -1142 463 -766
rect 497 -1142 513 -766
rect 447 -1154 513 -1142
rect 543 -766 605 -754
rect 543 -1142 559 -766
rect 593 -1142 605 -766
rect 543 -1154 605 -1142
<< pdiffc >>
rect -593 766 -559 1142
rect -497 766 -463 1142
rect -401 766 -367 1142
rect -305 766 -271 1142
rect -209 766 -175 1142
rect -113 766 -79 1142
rect -17 766 17 1142
rect 79 766 113 1142
rect 175 766 209 1142
rect 271 766 305 1142
rect 367 766 401 1142
rect 463 766 497 1142
rect 559 766 593 1142
rect -593 130 -559 506
rect -497 130 -463 506
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect 463 130 497 506
rect 559 130 593 506
rect -593 -506 -559 -130
rect -497 -506 -463 -130
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect 463 -506 497 -130
rect 559 -506 593 -130
rect -593 -1142 -559 -766
rect -497 -1142 -463 -766
rect -401 -1142 -367 -766
rect -305 -1142 -271 -766
rect -209 -1142 -175 -766
rect -113 -1142 -79 -766
rect -17 -1142 17 -766
rect 79 -1142 113 -766
rect 175 -1142 209 -766
rect 271 -1142 305 -766
rect 367 -1142 401 -766
rect 463 -1142 497 -766
rect 559 -1142 593 -766
<< nsubdiff >>
rect -707 1303 -611 1337
rect 611 1303 707 1337
rect -707 1241 -673 1303
rect 673 1241 707 1303
rect -707 -1303 -673 -1241
rect 673 -1303 707 -1241
rect -707 -1337 -611 -1303
rect 611 -1337 707 -1303
<< nsubdiffcont >>
rect -611 1303 611 1337
rect -707 -1241 -673 1241
rect 673 -1241 707 1241
rect -611 -1337 611 -1303
<< poly >>
rect -561 1235 -495 1251
rect -561 1201 -545 1235
rect -511 1201 -495 1235
rect -561 1185 -495 1201
rect -369 1235 -303 1251
rect -369 1201 -353 1235
rect -319 1201 -303 1235
rect -369 1185 -303 1201
rect -177 1235 -111 1251
rect -177 1201 -161 1235
rect -127 1201 -111 1235
rect -177 1185 -111 1201
rect 15 1235 81 1251
rect 15 1201 31 1235
rect 65 1201 81 1235
rect 15 1185 81 1201
rect 207 1235 273 1251
rect 207 1201 223 1235
rect 257 1201 273 1235
rect 207 1185 273 1201
rect 399 1235 465 1251
rect 399 1201 415 1235
rect 449 1201 465 1235
rect 399 1185 465 1201
rect -543 1154 -513 1185
rect -447 1154 -417 1180
rect -351 1154 -321 1185
rect -255 1154 -225 1180
rect -159 1154 -129 1185
rect -63 1154 -33 1180
rect 33 1154 63 1185
rect 129 1154 159 1180
rect 225 1154 255 1185
rect 321 1154 351 1180
rect 417 1154 447 1185
rect 513 1154 543 1180
rect -543 728 -513 754
rect -447 723 -417 754
rect -351 728 -321 754
rect -255 723 -225 754
rect -159 728 -129 754
rect -63 723 -33 754
rect 33 728 63 754
rect 129 723 159 754
rect 225 728 255 754
rect 321 723 351 754
rect 417 728 447 754
rect 513 723 543 754
rect -465 707 -399 723
rect -465 673 -449 707
rect -415 673 -399 707
rect -465 657 -399 673
rect -273 707 -207 723
rect -273 673 -257 707
rect -223 673 -207 707
rect -273 657 -207 673
rect -81 707 -15 723
rect -81 673 -65 707
rect -31 673 -15 707
rect -81 657 -15 673
rect 111 707 177 723
rect 111 673 127 707
rect 161 673 177 707
rect 111 657 177 673
rect 303 707 369 723
rect 303 673 319 707
rect 353 673 369 707
rect 303 657 369 673
rect 495 707 561 723
rect 495 673 511 707
rect 545 673 561 707
rect 495 657 561 673
rect -465 599 -399 615
rect -465 565 -449 599
rect -415 565 -399 599
rect -465 549 -399 565
rect -273 599 -207 615
rect -273 565 -257 599
rect -223 565 -207 599
rect -273 549 -207 565
rect -81 599 -15 615
rect -81 565 -65 599
rect -31 565 -15 599
rect -81 549 -15 565
rect 111 599 177 615
rect 111 565 127 599
rect 161 565 177 599
rect 111 549 177 565
rect 303 599 369 615
rect 303 565 319 599
rect 353 565 369 599
rect 303 549 369 565
rect 495 599 561 615
rect 495 565 511 599
rect 545 565 561 599
rect 495 549 561 565
rect -543 518 -513 544
rect -447 518 -417 549
rect -351 518 -321 544
rect -255 518 -225 549
rect -159 518 -129 544
rect -63 518 -33 549
rect 33 518 63 544
rect 129 518 159 549
rect 225 518 255 544
rect 321 518 351 549
rect 417 518 447 544
rect 513 518 543 549
rect -543 87 -513 118
rect -447 92 -417 118
rect -351 87 -321 118
rect -255 92 -225 118
rect -159 87 -129 118
rect -63 92 -33 118
rect 33 87 63 118
rect 129 92 159 118
rect 225 87 255 118
rect 321 92 351 118
rect 417 87 447 118
rect 513 92 543 118
rect -561 71 -495 87
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 399 -87 465 -71
rect -543 -118 -513 -87
rect -447 -118 -417 -92
rect -351 -118 -321 -87
rect -255 -118 -225 -92
rect -159 -118 -129 -87
rect -63 -118 -33 -92
rect 33 -118 63 -87
rect 129 -118 159 -92
rect 225 -118 255 -87
rect 321 -118 351 -92
rect 417 -118 447 -87
rect 513 -118 543 -92
rect -543 -544 -513 -518
rect -447 -549 -417 -518
rect -351 -544 -321 -518
rect -255 -549 -225 -518
rect -159 -544 -129 -518
rect -63 -549 -33 -518
rect 33 -544 63 -518
rect 129 -549 159 -518
rect 225 -544 255 -518
rect 321 -549 351 -518
rect 417 -544 447 -518
rect 513 -549 543 -518
rect -465 -565 -399 -549
rect -465 -599 -449 -565
rect -415 -599 -399 -565
rect -465 -615 -399 -599
rect -273 -565 -207 -549
rect -273 -599 -257 -565
rect -223 -599 -207 -565
rect -273 -615 -207 -599
rect -81 -565 -15 -549
rect -81 -599 -65 -565
rect -31 -599 -15 -565
rect -81 -615 -15 -599
rect 111 -565 177 -549
rect 111 -599 127 -565
rect 161 -599 177 -565
rect 111 -615 177 -599
rect 303 -565 369 -549
rect 303 -599 319 -565
rect 353 -599 369 -565
rect 303 -615 369 -599
rect 495 -565 561 -549
rect 495 -599 511 -565
rect 545 -599 561 -565
rect 495 -615 561 -599
rect -465 -673 -399 -657
rect -465 -707 -449 -673
rect -415 -707 -399 -673
rect -465 -723 -399 -707
rect -273 -673 -207 -657
rect -273 -707 -257 -673
rect -223 -707 -207 -673
rect -273 -723 -207 -707
rect -81 -673 -15 -657
rect -81 -707 -65 -673
rect -31 -707 -15 -673
rect -81 -723 -15 -707
rect 111 -673 177 -657
rect 111 -707 127 -673
rect 161 -707 177 -673
rect 111 -723 177 -707
rect 303 -673 369 -657
rect 303 -707 319 -673
rect 353 -707 369 -673
rect 303 -723 369 -707
rect 495 -673 561 -657
rect 495 -707 511 -673
rect 545 -707 561 -673
rect 495 -723 561 -707
rect -543 -754 -513 -728
rect -447 -754 -417 -723
rect -351 -754 -321 -728
rect -255 -754 -225 -723
rect -159 -754 -129 -728
rect -63 -754 -33 -723
rect 33 -754 63 -728
rect 129 -754 159 -723
rect 225 -754 255 -728
rect 321 -754 351 -723
rect 417 -754 447 -728
rect 513 -754 543 -723
rect -543 -1185 -513 -1154
rect -447 -1180 -417 -1154
rect -351 -1185 -321 -1154
rect -255 -1180 -225 -1154
rect -159 -1185 -129 -1154
rect -63 -1180 -33 -1154
rect 33 -1185 63 -1154
rect 129 -1180 159 -1154
rect 225 -1185 255 -1154
rect 321 -1180 351 -1154
rect 417 -1185 447 -1154
rect 513 -1180 543 -1154
rect -561 -1201 -495 -1185
rect -561 -1235 -545 -1201
rect -511 -1235 -495 -1201
rect -561 -1251 -495 -1235
rect -369 -1201 -303 -1185
rect -369 -1235 -353 -1201
rect -319 -1235 -303 -1201
rect -369 -1251 -303 -1235
rect -177 -1201 -111 -1185
rect -177 -1235 -161 -1201
rect -127 -1235 -111 -1201
rect -177 -1251 -111 -1235
rect 15 -1201 81 -1185
rect 15 -1235 31 -1201
rect 65 -1235 81 -1201
rect 15 -1251 81 -1235
rect 207 -1201 273 -1185
rect 207 -1235 223 -1201
rect 257 -1235 273 -1201
rect 207 -1251 273 -1235
rect 399 -1201 465 -1185
rect 399 -1235 415 -1201
rect 449 -1235 465 -1201
rect 399 -1251 465 -1235
<< polycont >>
rect -545 1201 -511 1235
rect -353 1201 -319 1235
rect -161 1201 -127 1235
rect 31 1201 65 1235
rect 223 1201 257 1235
rect 415 1201 449 1235
rect -449 673 -415 707
rect -257 673 -223 707
rect -65 673 -31 707
rect 127 673 161 707
rect 319 673 353 707
rect 511 673 545 707
rect -449 565 -415 599
rect -257 565 -223 599
rect -65 565 -31 599
rect 127 565 161 599
rect 319 565 353 599
rect 511 565 545 599
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -449 -599 -415 -565
rect -257 -599 -223 -565
rect -65 -599 -31 -565
rect 127 -599 161 -565
rect 319 -599 353 -565
rect 511 -599 545 -565
rect -449 -707 -415 -673
rect -257 -707 -223 -673
rect -65 -707 -31 -673
rect 127 -707 161 -673
rect 319 -707 353 -673
rect 511 -707 545 -673
rect -545 -1235 -511 -1201
rect -353 -1235 -319 -1201
rect -161 -1235 -127 -1201
rect 31 -1235 65 -1201
rect 223 -1235 257 -1201
rect 415 -1235 449 -1201
<< locali >>
rect -707 1303 -611 1337
rect 611 1303 707 1337
rect -707 1241 -673 1303
rect 673 1241 707 1303
rect -561 1201 -545 1235
rect -511 1201 -495 1235
rect -369 1201 -353 1235
rect -319 1201 -303 1235
rect -177 1201 -161 1235
rect -127 1201 -111 1235
rect 15 1201 31 1235
rect 65 1201 81 1235
rect 207 1201 223 1235
rect 257 1201 273 1235
rect 399 1201 415 1235
rect 449 1201 465 1235
rect -593 1142 -559 1158
rect -593 750 -559 766
rect -497 1142 -463 1158
rect -497 750 -463 766
rect -401 1142 -367 1158
rect -401 750 -367 766
rect -305 1142 -271 1158
rect -305 750 -271 766
rect -209 1142 -175 1158
rect -209 750 -175 766
rect -113 1142 -79 1158
rect -113 750 -79 766
rect -17 1142 17 1158
rect -17 750 17 766
rect 79 1142 113 1158
rect 79 750 113 766
rect 175 1142 209 1158
rect 175 750 209 766
rect 271 1142 305 1158
rect 271 750 305 766
rect 367 1142 401 1158
rect 367 750 401 766
rect 463 1142 497 1158
rect 463 750 497 766
rect 559 1142 593 1158
rect 559 750 593 766
rect -465 673 -449 707
rect -415 673 -399 707
rect -273 673 -257 707
rect -223 673 -207 707
rect -81 673 -65 707
rect -31 673 -15 707
rect 111 673 127 707
rect 161 673 177 707
rect 303 673 319 707
rect 353 673 369 707
rect 495 673 511 707
rect 545 673 561 707
rect -465 565 -449 599
rect -415 565 -399 599
rect -273 565 -257 599
rect -223 565 -207 599
rect -81 565 -65 599
rect -31 565 -15 599
rect 111 565 127 599
rect 161 565 177 599
rect 303 565 319 599
rect 353 565 369 599
rect 495 565 511 599
rect 545 565 561 599
rect -593 506 -559 522
rect -593 114 -559 130
rect -497 506 -463 522
rect -497 114 -463 130
rect -401 506 -367 522
rect -401 114 -367 130
rect -305 506 -271 522
rect -305 114 -271 130
rect -209 506 -175 522
rect -209 114 -175 130
rect -113 506 -79 522
rect -113 114 -79 130
rect -17 506 17 522
rect -17 114 17 130
rect 79 506 113 522
rect 79 114 113 130
rect 175 506 209 522
rect 175 114 209 130
rect 271 506 305 522
rect 271 114 305 130
rect 367 506 401 522
rect 367 114 401 130
rect 463 506 497 522
rect 463 114 497 130
rect 559 506 593 522
rect 559 114 593 130
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect -593 -130 -559 -114
rect -593 -522 -559 -506
rect -497 -130 -463 -114
rect -497 -522 -463 -506
rect -401 -130 -367 -114
rect -401 -522 -367 -506
rect -305 -130 -271 -114
rect -305 -522 -271 -506
rect -209 -130 -175 -114
rect -209 -522 -175 -506
rect -113 -130 -79 -114
rect -113 -522 -79 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 79 -130 113 -114
rect 79 -522 113 -506
rect 175 -130 209 -114
rect 175 -522 209 -506
rect 271 -130 305 -114
rect 271 -522 305 -506
rect 367 -130 401 -114
rect 367 -522 401 -506
rect 463 -130 497 -114
rect 463 -522 497 -506
rect 559 -130 593 -114
rect 559 -522 593 -506
rect -465 -599 -449 -565
rect -415 -599 -399 -565
rect -273 -599 -257 -565
rect -223 -599 -207 -565
rect -81 -599 -65 -565
rect -31 -599 -15 -565
rect 111 -599 127 -565
rect 161 -599 177 -565
rect 303 -599 319 -565
rect 353 -599 369 -565
rect 495 -599 511 -565
rect 545 -599 561 -565
rect -465 -707 -449 -673
rect -415 -707 -399 -673
rect -273 -707 -257 -673
rect -223 -707 -207 -673
rect -81 -707 -65 -673
rect -31 -707 -15 -673
rect 111 -707 127 -673
rect 161 -707 177 -673
rect 303 -707 319 -673
rect 353 -707 369 -673
rect 495 -707 511 -673
rect 545 -707 561 -673
rect -593 -766 -559 -750
rect -593 -1158 -559 -1142
rect -497 -766 -463 -750
rect -497 -1158 -463 -1142
rect -401 -766 -367 -750
rect -401 -1158 -367 -1142
rect -305 -766 -271 -750
rect -305 -1158 -271 -1142
rect -209 -766 -175 -750
rect -209 -1158 -175 -1142
rect -113 -766 -79 -750
rect -113 -1158 -79 -1142
rect -17 -766 17 -750
rect -17 -1158 17 -1142
rect 79 -766 113 -750
rect 79 -1158 113 -1142
rect 175 -766 209 -750
rect 175 -1158 209 -1142
rect 271 -766 305 -750
rect 271 -1158 305 -1142
rect 367 -766 401 -750
rect 367 -1158 401 -1142
rect 463 -766 497 -750
rect 463 -1158 497 -1142
rect 559 -766 593 -750
rect 559 -1158 593 -1142
rect -561 -1235 -545 -1201
rect -511 -1235 -495 -1201
rect -369 -1235 -353 -1201
rect -319 -1235 -303 -1201
rect -177 -1235 -161 -1201
rect -127 -1235 -111 -1201
rect 15 -1235 31 -1201
rect 65 -1235 81 -1201
rect 207 -1235 223 -1201
rect 257 -1235 273 -1201
rect 399 -1235 415 -1201
rect 449 -1235 465 -1201
rect -707 -1303 -673 -1241
rect 673 -1303 707 -1241
rect -707 -1337 -611 -1303
rect 611 -1337 707 -1303
<< viali >>
rect -545 1201 -511 1235
rect -353 1201 -319 1235
rect -161 1201 -127 1235
rect 31 1201 65 1235
rect 223 1201 257 1235
rect 415 1201 449 1235
rect -593 766 -559 1142
rect -497 766 -463 1142
rect -401 766 -367 1142
rect -305 766 -271 1142
rect -209 766 -175 1142
rect -113 766 -79 1142
rect -17 766 17 1142
rect 79 766 113 1142
rect 175 766 209 1142
rect 271 766 305 1142
rect 367 766 401 1142
rect 463 766 497 1142
rect 559 766 593 1142
rect -449 673 -415 707
rect -257 673 -223 707
rect -65 673 -31 707
rect 127 673 161 707
rect 319 673 353 707
rect 511 673 545 707
rect -449 565 -415 599
rect -257 565 -223 599
rect -65 565 -31 599
rect 127 565 161 599
rect 319 565 353 599
rect 511 565 545 599
rect -593 130 -559 506
rect -497 130 -463 506
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect 463 130 497 506
rect 559 130 593 506
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -593 -506 -559 -130
rect -497 -506 -463 -130
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect 463 -506 497 -130
rect 559 -506 593 -130
rect -449 -599 -415 -565
rect -257 -599 -223 -565
rect -65 -599 -31 -565
rect 127 -599 161 -565
rect 319 -599 353 -565
rect 511 -599 545 -565
rect -449 -707 -415 -673
rect -257 -707 -223 -673
rect -65 -707 -31 -673
rect 127 -707 161 -673
rect 319 -707 353 -673
rect 511 -707 545 -673
rect -593 -1142 -559 -766
rect -497 -1142 -463 -766
rect -401 -1142 -367 -766
rect -305 -1142 -271 -766
rect -209 -1142 -175 -766
rect -113 -1142 -79 -766
rect -17 -1142 17 -766
rect 79 -1142 113 -766
rect 175 -1142 209 -766
rect 271 -1142 305 -766
rect 367 -1142 401 -766
rect 463 -1142 497 -766
rect 559 -1142 593 -766
rect -545 -1235 -511 -1201
rect -353 -1235 -319 -1201
rect -161 -1235 -127 -1201
rect 31 -1235 65 -1201
rect 223 -1235 257 -1201
rect 415 -1235 449 -1201
<< metal1 >>
rect -557 1235 -499 1241
rect -557 1201 -545 1235
rect -511 1201 -499 1235
rect -557 1195 -499 1201
rect -365 1235 -307 1241
rect -365 1201 -353 1235
rect -319 1201 -307 1235
rect -365 1195 -307 1201
rect -173 1235 -115 1241
rect -173 1201 -161 1235
rect -127 1201 -115 1235
rect -173 1195 -115 1201
rect 19 1235 77 1241
rect 19 1201 31 1235
rect 65 1201 77 1235
rect 19 1195 77 1201
rect 211 1235 269 1241
rect 211 1201 223 1235
rect 257 1201 269 1235
rect 211 1195 269 1201
rect 403 1235 461 1241
rect 403 1201 415 1235
rect 449 1201 461 1235
rect 403 1195 461 1201
rect -599 1142 -553 1154
rect -599 766 -593 1142
rect -559 766 -553 1142
rect -599 754 -553 766
rect -503 1142 -457 1154
rect -503 766 -497 1142
rect -463 766 -457 1142
rect -503 754 -457 766
rect -407 1142 -361 1154
rect -407 766 -401 1142
rect -367 766 -361 1142
rect -407 754 -361 766
rect -311 1142 -265 1154
rect -311 766 -305 1142
rect -271 766 -265 1142
rect -311 754 -265 766
rect -215 1142 -169 1154
rect -215 766 -209 1142
rect -175 766 -169 1142
rect -215 754 -169 766
rect -119 1142 -73 1154
rect -119 766 -113 1142
rect -79 766 -73 1142
rect -119 754 -73 766
rect -23 1142 23 1154
rect -23 766 -17 1142
rect 17 766 23 1142
rect -23 754 23 766
rect 73 1142 119 1154
rect 73 766 79 1142
rect 113 766 119 1142
rect 73 754 119 766
rect 169 1142 215 1154
rect 169 766 175 1142
rect 209 766 215 1142
rect 169 754 215 766
rect 265 1142 311 1154
rect 265 766 271 1142
rect 305 766 311 1142
rect 265 754 311 766
rect 361 1142 407 1154
rect 361 766 367 1142
rect 401 766 407 1142
rect 361 754 407 766
rect 457 1142 503 1154
rect 457 766 463 1142
rect 497 766 503 1142
rect 457 754 503 766
rect 553 1142 599 1154
rect 553 766 559 1142
rect 593 766 599 1142
rect 553 754 599 766
rect -461 707 -403 713
rect -461 673 -449 707
rect -415 673 -403 707
rect -461 667 -403 673
rect -269 707 -211 713
rect -269 673 -257 707
rect -223 673 -211 707
rect -269 667 -211 673
rect -77 707 -19 713
rect -77 673 -65 707
rect -31 673 -19 707
rect -77 667 -19 673
rect 115 707 173 713
rect 115 673 127 707
rect 161 673 173 707
rect 115 667 173 673
rect 307 707 365 713
rect 307 673 319 707
rect 353 673 365 707
rect 307 667 365 673
rect 499 707 557 713
rect 499 673 511 707
rect 545 673 557 707
rect 499 667 557 673
rect -461 599 -403 605
rect -461 565 -449 599
rect -415 565 -403 599
rect -461 559 -403 565
rect -269 599 -211 605
rect -269 565 -257 599
rect -223 565 -211 599
rect -269 559 -211 565
rect -77 599 -19 605
rect -77 565 -65 599
rect -31 565 -19 599
rect -77 559 -19 565
rect 115 599 173 605
rect 115 565 127 599
rect 161 565 173 599
rect 115 559 173 565
rect 307 599 365 605
rect 307 565 319 599
rect 353 565 365 599
rect 307 559 365 565
rect 499 599 557 605
rect 499 565 511 599
rect 545 565 557 599
rect 499 559 557 565
rect -599 506 -553 518
rect -599 130 -593 506
rect -559 130 -553 506
rect -599 118 -553 130
rect -503 506 -457 518
rect -503 130 -497 506
rect -463 130 -457 506
rect -503 118 -457 130
rect -407 506 -361 518
rect -407 130 -401 506
rect -367 130 -361 506
rect -407 118 -361 130
rect -311 506 -265 518
rect -311 130 -305 506
rect -271 130 -265 506
rect -311 118 -265 130
rect -215 506 -169 518
rect -215 130 -209 506
rect -175 130 -169 506
rect -215 118 -169 130
rect -119 506 -73 518
rect -119 130 -113 506
rect -79 130 -73 506
rect -119 118 -73 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 73 506 119 518
rect 73 130 79 506
rect 113 130 119 506
rect 73 118 119 130
rect 169 506 215 518
rect 169 130 175 506
rect 209 130 215 506
rect 169 118 215 130
rect 265 506 311 518
rect 265 130 271 506
rect 305 130 311 506
rect 265 118 311 130
rect 361 506 407 518
rect 361 130 367 506
rect 401 130 407 506
rect 361 118 407 130
rect 457 506 503 518
rect 457 130 463 506
rect 497 130 503 506
rect 457 118 503 130
rect 553 506 599 518
rect 553 130 559 506
rect 593 130 599 506
rect 553 118 599 130
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect -599 -130 -553 -118
rect -599 -506 -593 -130
rect -559 -506 -553 -130
rect -599 -518 -553 -506
rect -503 -130 -457 -118
rect -503 -506 -497 -130
rect -463 -506 -457 -130
rect -503 -518 -457 -506
rect -407 -130 -361 -118
rect -407 -506 -401 -130
rect -367 -506 -361 -130
rect -407 -518 -361 -506
rect -311 -130 -265 -118
rect -311 -506 -305 -130
rect -271 -506 -265 -130
rect -311 -518 -265 -506
rect -215 -130 -169 -118
rect -215 -506 -209 -130
rect -175 -506 -169 -130
rect -215 -518 -169 -506
rect -119 -130 -73 -118
rect -119 -506 -113 -130
rect -79 -506 -73 -130
rect -119 -518 -73 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 73 -130 119 -118
rect 73 -506 79 -130
rect 113 -506 119 -130
rect 73 -518 119 -506
rect 169 -130 215 -118
rect 169 -506 175 -130
rect 209 -506 215 -130
rect 169 -518 215 -506
rect 265 -130 311 -118
rect 265 -506 271 -130
rect 305 -506 311 -130
rect 265 -518 311 -506
rect 361 -130 407 -118
rect 361 -506 367 -130
rect 401 -506 407 -130
rect 361 -518 407 -506
rect 457 -130 503 -118
rect 457 -506 463 -130
rect 497 -506 503 -130
rect 457 -518 503 -506
rect 553 -130 599 -118
rect 553 -506 559 -130
rect 593 -506 599 -130
rect 553 -518 599 -506
rect -461 -565 -403 -559
rect -461 -599 -449 -565
rect -415 -599 -403 -565
rect -461 -605 -403 -599
rect -269 -565 -211 -559
rect -269 -599 -257 -565
rect -223 -599 -211 -565
rect -269 -605 -211 -599
rect -77 -565 -19 -559
rect -77 -599 -65 -565
rect -31 -599 -19 -565
rect -77 -605 -19 -599
rect 115 -565 173 -559
rect 115 -599 127 -565
rect 161 -599 173 -565
rect 115 -605 173 -599
rect 307 -565 365 -559
rect 307 -599 319 -565
rect 353 -599 365 -565
rect 307 -605 365 -599
rect 499 -565 557 -559
rect 499 -599 511 -565
rect 545 -599 557 -565
rect 499 -605 557 -599
rect -461 -673 -403 -667
rect -461 -707 -449 -673
rect -415 -707 -403 -673
rect -461 -713 -403 -707
rect -269 -673 -211 -667
rect -269 -707 -257 -673
rect -223 -707 -211 -673
rect -269 -713 -211 -707
rect -77 -673 -19 -667
rect -77 -707 -65 -673
rect -31 -707 -19 -673
rect -77 -713 -19 -707
rect 115 -673 173 -667
rect 115 -707 127 -673
rect 161 -707 173 -673
rect 115 -713 173 -707
rect 307 -673 365 -667
rect 307 -707 319 -673
rect 353 -707 365 -673
rect 307 -713 365 -707
rect 499 -673 557 -667
rect 499 -707 511 -673
rect 545 -707 557 -673
rect 499 -713 557 -707
rect -599 -766 -553 -754
rect -599 -1142 -593 -766
rect -559 -1142 -553 -766
rect -599 -1154 -553 -1142
rect -503 -766 -457 -754
rect -503 -1142 -497 -766
rect -463 -1142 -457 -766
rect -503 -1154 -457 -1142
rect -407 -766 -361 -754
rect -407 -1142 -401 -766
rect -367 -1142 -361 -766
rect -407 -1154 -361 -1142
rect -311 -766 -265 -754
rect -311 -1142 -305 -766
rect -271 -1142 -265 -766
rect -311 -1154 -265 -1142
rect -215 -766 -169 -754
rect -215 -1142 -209 -766
rect -175 -1142 -169 -766
rect -215 -1154 -169 -1142
rect -119 -766 -73 -754
rect -119 -1142 -113 -766
rect -79 -1142 -73 -766
rect -119 -1154 -73 -1142
rect -23 -766 23 -754
rect -23 -1142 -17 -766
rect 17 -1142 23 -766
rect -23 -1154 23 -1142
rect 73 -766 119 -754
rect 73 -1142 79 -766
rect 113 -1142 119 -766
rect 73 -1154 119 -1142
rect 169 -766 215 -754
rect 169 -1142 175 -766
rect 209 -1142 215 -766
rect 169 -1154 215 -1142
rect 265 -766 311 -754
rect 265 -1142 271 -766
rect 305 -1142 311 -766
rect 265 -1154 311 -1142
rect 361 -766 407 -754
rect 361 -1142 367 -766
rect 401 -1142 407 -766
rect 361 -1154 407 -1142
rect 457 -766 503 -754
rect 457 -1142 463 -766
rect 497 -1142 503 -766
rect 457 -1154 503 -1142
rect 553 -766 599 -754
rect 553 -1142 559 -766
rect 593 -1142 599 -766
rect 553 -1154 599 -1142
rect -557 -1201 -499 -1195
rect -557 -1235 -545 -1201
rect -511 -1235 -499 -1201
rect -557 -1241 -499 -1235
rect -365 -1201 -307 -1195
rect -365 -1235 -353 -1201
rect -319 -1235 -307 -1201
rect -365 -1241 -307 -1235
rect -173 -1201 -115 -1195
rect -173 -1235 -161 -1201
rect -127 -1235 -115 -1201
rect -173 -1241 -115 -1235
rect 19 -1201 77 -1195
rect 19 -1235 31 -1201
rect 65 -1235 77 -1201
rect 19 -1241 77 -1235
rect 211 -1201 269 -1195
rect 211 -1235 223 -1201
rect 257 -1235 269 -1201
rect 211 -1241 269 -1235
rect 403 -1201 461 -1195
rect 403 -1235 415 -1201
rect 449 -1235 461 -1201
rect 403 -1241 461 -1235
<< properties >>
string FIXED_BBOX -690 -1320 690 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 4 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
