magic
tech sky130A
magscale 1 2
timestamp 1645790779
<< error_p >>
rect -2381 1199 -2323 1205
rect -2189 1199 -2131 1205
rect -1997 1199 -1939 1205
rect -1805 1199 -1747 1205
rect -1613 1199 -1555 1205
rect -1421 1199 -1363 1205
rect -1229 1199 -1171 1205
rect -1037 1199 -979 1205
rect -845 1199 -787 1205
rect -653 1199 -595 1205
rect -461 1199 -403 1205
rect -269 1199 -211 1205
rect -77 1199 -19 1205
rect 115 1199 173 1205
rect 307 1199 365 1205
rect 499 1199 557 1205
rect 691 1199 749 1205
rect 883 1199 941 1205
rect 1075 1199 1133 1205
rect 1267 1199 1325 1205
rect 1459 1199 1517 1205
rect 1651 1199 1709 1205
rect 1843 1199 1901 1205
rect 2035 1199 2093 1205
rect 2227 1199 2285 1205
rect -2381 1165 -2369 1199
rect -2189 1165 -2177 1199
rect -1997 1165 -1985 1199
rect -1805 1165 -1793 1199
rect -1613 1165 -1601 1199
rect -1421 1165 -1409 1199
rect -1229 1165 -1217 1199
rect -1037 1165 -1025 1199
rect -845 1165 -833 1199
rect -653 1165 -641 1199
rect -461 1165 -449 1199
rect -269 1165 -257 1199
rect -77 1165 -65 1199
rect 115 1165 127 1199
rect 307 1165 319 1199
rect 499 1165 511 1199
rect 691 1165 703 1199
rect 883 1165 895 1199
rect 1075 1165 1087 1199
rect 1267 1165 1279 1199
rect 1459 1165 1471 1199
rect 1651 1165 1663 1199
rect 1843 1165 1855 1199
rect 2035 1165 2047 1199
rect 2227 1165 2239 1199
rect -2381 1159 -2323 1165
rect -2189 1159 -2131 1165
rect -1997 1159 -1939 1165
rect -1805 1159 -1747 1165
rect -1613 1159 -1555 1165
rect -1421 1159 -1363 1165
rect -1229 1159 -1171 1165
rect -1037 1159 -979 1165
rect -845 1159 -787 1165
rect -653 1159 -595 1165
rect -461 1159 -403 1165
rect -269 1159 -211 1165
rect -77 1159 -19 1165
rect 115 1159 173 1165
rect 307 1159 365 1165
rect 499 1159 557 1165
rect 691 1159 749 1165
rect 883 1159 941 1165
rect 1075 1159 1133 1165
rect 1267 1159 1325 1165
rect 1459 1159 1517 1165
rect 1651 1159 1709 1165
rect 1843 1159 1901 1165
rect 2035 1159 2093 1165
rect 2227 1159 2285 1165
rect -2285 689 -2227 695
rect -2093 689 -2035 695
rect -1901 689 -1843 695
rect -1709 689 -1651 695
rect -1517 689 -1459 695
rect -1325 689 -1267 695
rect -1133 689 -1075 695
rect -941 689 -883 695
rect -749 689 -691 695
rect -557 689 -499 695
rect -365 689 -307 695
rect -173 689 -115 695
rect 19 689 77 695
rect 211 689 269 695
rect 403 689 461 695
rect 595 689 653 695
rect 787 689 845 695
rect 979 689 1037 695
rect 1171 689 1229 695
rect 1363 689 1421 695
rect 1555 689 1613 695
rect 1747 689 1805 695
rect 1939 689 1997 695
rect 2131 689 2189 695
rect 2323 689 2381 695
rect -2285 655 -2273 689
rect -2093 655 -2081 689
rect -1901 655 -1889 689
rect -1709 655 -1697 689
rect -1517 655 -1505 689
rect -1325 655 -1313 689
rect -1133 655 -1121 689
rect -941 655 -929 689
rect -749 655 -737 689
rect -557 655 -545 689
rect -365 655 -353 689
rect -173 655 -161 689
rect 19 655 31 689
rect 211 655 223 689
rect 403 655 415 689
rect 595 655 607 689
rect 787 655 799 689
rect 979 655 991 689
rect 1171 655 1183 689
rect 1363 655 1375 689
rect 1555 655 1567 689
rect 1747 655 1759 689
rect 1939 655 1951 689
rect 2131 655 2143 689
rect 2323 655 2335 689
rect -2285 649 -2227 655
rect -2093 649 -2035 655
rect -1901 649 -1843 655
rect -1709 649 -1651 655
rect -1517 649 -1459 655
rect -1325 649 -1267 655
rect -1133 649 -1075 655
rect -941 649 -883 655
rect -749 649 -691 655
rect -557 649 -499 655
rect -365 649 -307 655
rect -173 649 -115 655
rect 19 649 77 655
rect 211 649 269 655
rect 403 649 461 655
rect 595 649 653 655
rect 787 649 845 655
rect 979 649 1037 655
rect 1171 649 1229 655
rect 1363 649 1421 655
rect 1555 649 1613 655
rect 1747 649 1805 655
rect 1939 649 1997 655
rect 2131 649 2189 655
rect 2323 649 2381 655
rect -2285 581 -2227 587
rect -2093 581 -2035 587
rect -1901 581 -1843 587
rect -1709 581 -1651 587
rect -1517 581 -1459 587
rect -1325 581 -1267 587
rect -1133 581 -1075 587
rect -941 581 -883 587
rect -749 581 -691 587
rect -557 581 -499 587
rect -365 581 -307 587
rect -173 581 -115 587
rect 19 581 77 587
rect 211 581 269 587
rect 403 581 461 587
rect 595 581 653 587
rect 787 581 845 587
rect 979 581 1037 587
rect 1171 581 1229 587
rect 1363 581 1421 587
rect 1555 581 1613 587
rect 1747 581 1805 587
rect 1939 581 1997 587
rect 2131 581 2189 587
rect 2323 581 2381 587
rect -2285 547 -2273 581
rect -2093 547 -2081 581
rect -1901 547 -1889 581
rect -1709 547 -1697 581
rect -1517 547 -1505 581
rect -1325 547 -1313 581
rect -1133 547 -1121 581
rect -941 547 -929 581
rect -749 547 -737 581
rect -557 547 -545 581
rect -365 547 -353 581
rect -173 547 -161 581
rect 19 547 31 581
rect 211 547 223 581
rect 403 547 415 581
rect 595 547 607 581
rect 787 547 799 581
rect 979 547 991 581
rect 1171 547 1183 581
rect 1363 547 1375 581
rect 1555 547 1567 581
rect 1747 547 1759 581
rect 1939 547 1951 581
rect 2131 547 2143 581
rect 2323 547 2335 581
rect -2285 541 -2227 547
rect -2093 541 -2035 547
rect -1901 541 -1843 547
rect -1709 541 -1651 547
rect -1517 541 -1459 547
rect -1325 541 -1267 547
rect -1133 541 -1075 547
rect -941 541 -883 547
rect -749 541 -691 547
rect -557 541 -499 547
rect -365 541 -307 547
rect -173 541 -115 547
rect 19 541 77 547
rect 211 541 269 547
rect 403 541 461 547
rect 595 541 653 547
rect 787 541 845 547
rect 979 541 1037 547
rect 1171 541 1229 547
rect 1363 541 1421 547
rect 1555 541 1613 547
rect 1747 541 1805 547
rect 1939 541 1997 547
rect 2131 541 2189 547
rect 2323 541 2381 547
rect -2381 71 -2323 77
rect -2189 71 -2131 77
rect -1997 71 -1939 77
rect -1805 71 -1747 77
rect -1613 71 -1555 77
rect -1421 71 -1363 77
rect -1229 71 -1171 77
rect -1037 71 -979 77
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect 1075 71 1133 77
rect 1267 71 1325 77
rect 1459 71 1517 77
rect 1651 71 1709 77
rect 1843 71 1901 77
rect 2035 71 2093 77
rect 2227 71 2285 77
rect -2381 37 -2369 71
rect -2189 37 -2177 71
rect -1997 37 -1985 71
rect -1805 37 -1793 71
rect -1613 37 -1601 71
rect -1421 37 -1409 71
rect -1229 37 -1217 71
rect -1037 37 -1025 71
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect 1075 37 1087 71
rect 1267 37 1279 71
rect 1459 37 1471 71
rect 1651 37 1663 71
rect 1843 37 1855 71
rect 2035 37 2047 71
rect 2227 37 2239 71
rect -2381 31 -2323 37
rect -2189 31 -2131 37
rect -1997 31 -1939 37
rect -1805 31 -1747 37
rect -1613 31 -1555 37
rect -1421 31 -1363 37
rect -1229 31 -1171 37
rect -1037 31 -979 37
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect 1075 31 1133 37
rect 1267 31 1325 37
rect 1459 31 1517 37
rect 1651 31 1709 37
rect 1843 31 1901 37
rect 2035 31 2093 37
rect 2227 31 2285 37
rect -2381 -37 -2323 -31
rect -2189 -37 -2131 -31
rect -1997 -37 -1939 -31
rect -1805 -37 -1747 -31
rect -1613 -37 -1555 -31
rect -1421 -37 -1363 -31
rect -1229 -37 -1171 -31
rect -1037 -37 -979 -31
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect 1075 -37 1133 -31
rect 1267 -37 1325 -31
rect 1459 -37 1517 -31
rect 1651 -37 1709 -31
rect 1843 -37 1901 -31
rect 2035 -37 2093 -31
rect 2227 -37 2285 -31
rect -2381 -71 -2369 -37
rect -2189 -71 -2177 -37
rect -1997 -71 -1985 -37
rect -1805 -71 -1793 -37
rect -1613 -71 -1601 -37
rect -1421 -71 -1409 -37
rect -1229 -71 -1217 -37
rect -1037 -71 -1025 -37
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect 1075 -71 1087 -37
rect 1267 -71 1279 -37
rect 1459 -71 1471 -37
rect 1651 -71 1663 -37
rect 1843 -71 1855 -37
rect 2035 -71 2047 -37
rect 2227 -71 2239 -37
rect -2381 -77 -2323 -71
rect -2189 -77 -2131 -71
rect -1997 -77 -1939 -71
rect -1805 -77 -1747 -71
rect -1613 -77 -1555 -71
rect -1421 -77 -1363 -71
rect -1229 -77 -1171 -71
rect -1037 -77 -979 -71
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect 1075 -77 1133 -71
rect 1267 -77 1325 -71
rect 1459 -77 1517 -71
rect 1651 -77 1709 -71
rect 1843 -77 1901 -71
rect 2035 -77 2093 -71
rect 2227 -77 2285 -71
rect -2285 -547 -2227 -541
rect -2093 -547 -2035 -541
rect -1901 -547 -1843 -541
rect -1709 -547 -1651 -541
rect -1517 -547 -1459 -541
rect -1325 -547 -1267 -541
rect -1133 -547 -1075 -541
rect -941 -547 -883 -541
rect -749 -547 -691 -541
rect -557 -547 -499 -541
rect -365 -547 -307 -541
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect 211 -547 269 -541
rect 403 -547 461 -541
rect 595 -547 653 -541
rect 787 -547 845 -541
rect 979 -547 1037 -541
rect 1171 -547 1229 -541
rect 1363 -547 1421 -541
rect 1555 -547 1613 -541
rect 1747 -547 1805 -541
rect 1939 -547 1997 -541
rect 2131 -547 2189 -541
rect 2323 -547 2381 -541
rect -2285 -581 -2273 -547
rect -2093 -581 -2081 -547
rect -1901 -581 -1889 -547
rect -1709 -581 -1697 -547
rect -1517 -581 -1505 -547
rect -1325 -581 -1313 -547
rect -1133 -581 -1121 -547
rect -941 -581 -929 -547
rect -749 -581 -737 -547
rect -557 -581 -545 -547
rect -365 -581 -353 -547
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect 211 -581 223 -547
rect 403 -581 415 -547
rect 595 -581 607 -547
rect 787 -581 799 -547
rect 979 -581 991 -547
rect 1171 -581 1183 -547
rect 1363 -581 1375 -547
rect 1555 -581 1567 -547
rect 1747 -581 1759 -547
rect 1939 -581 1951 -547
rect 2131 -581 2143 -547
rect 2323 -581 2335 -547
rect -2285 -587 -2227 -581
rect -2093 -587 -2035 -581
rect -1901 -587 -1843 -581
rect -1709 -587 -1651 -581
rect -1517 -587 -1459 -581
rect -1325 -587 -1267 -581
rect -1133 -587 -1075 -581
rect -941 -587 -883 -581
rect -749 -587 -691 -581
rect -557 -587 -499 -581
rect -365 -587 -307 -581
rect -173 -587 -115 -581
rect 19 -587 77 -581
rect 211 -587 269 -581
rect 403 -587 461 -581
rect 595 -587 653 -581
rect 787 -587 845 -581
rect 979 -587 1037 -581
rect 1171 -587 1229 -581
rect 1363 -587 1421 -581
rect 1555 -587 1613 -581
rect 1747 -587 1805 -581
rect 1939 -587 1997 -581
rect 2131 -587 2189 -581
rect 2323 -587 2381 -581
rect -2285 -655 -2227 -649
rect -2093 -655 -2035 -649
rect -1901 -655 -1843 -649
rect -1709 -655 -1651 -649
rect -1517 -655 -1459 -649
rect -1325 -655 -1267 -649
rect -1133 -655 -1075 -649
rect -941 -655 -883 -649
rect -749 -655 -691 -649
rect -557 -655 -499 -649
rect -365 -655 -307 -649
rect -173 -655 -115 -649
rect 19 -655 77 -649
rect 211 -655 269 -649
rect 403 -655 461 -649
rect 595 -655 653 -649
rect 787 -655 845 -649
rect 979 -655 1037 -649
rect 1171 -655 1229 -649
rect 1363 -655 1421 -649
rect 1555 -655 1613 -649
rect 1747 -655 1805 -649
rect 1939 -655 1997 -649
rect 2131 -655 2189 -649
rect 2323 -655 2381 -649
rect -2285 -689 -2273 -655
rect -2093 -689 -2081 -655
rect -1901 -689 -1889 -655
rect -1709 -689 -1697 -655
rect -1517 -689 -1505 -655
rect -1325 -689 -1313 -655
rect -1133 -689 -1121 -655
rect -941 -689 -929 -655
rect -749 -689 -737 -655
rect -557 -689 -545 -655
rect -365 -689 -353 -655
rect -173 -689 -161 -655
rect 19 -689 31 -655
rect 211 -689 223 -655
rect 403 -689 415 -655
rect 595 -689 607 -655
rect 787 -689 799 -655
rect 979 -689 991 -655
rect 1171 -689 1183 -655
rect 1363 -689 1375 -655
rect 1555 -689 1567 -655
rect 1747 -689 1759 -655
rect 1939 -689 1951 -655
rect 2131 -689 2143 -655
rect 2323 -689 2335 -655
rect -2285 -695 -2227 -689
rect -2093 -695 -2035 -689
rect -1901 -695 -1843 -689
rect -1709 -695 -1651 -689
rect -1517 -695 -1459 -689
rect -1325 -695 -1267 -689
rect -1133 -695 -1075 -689
rect -941 -695 -883 -689
rect -749 -695 -691 -689
rect -557 -695 -499 -689
rect -365 -695 -307 -689
rect -173 -695 -115 -689
rect 19 -695 77 -689
rect 211 -695 269 -689
rect 403 -695 461 -689
rect 595 -695 653 -689
rect 787 -695 845 -689
rect 979 -695 1037 -689
rect 1171 -695 1229 -689
rect 1363 -695 1421 -689
rect 1555 -695 1613 -689
rect 1747 -695 1805 -689
rect 1939 -695 1997 -689
rect 2131 -695 2189 -689
rect 2323 -695 2381 -689
rect -2381 -1165 -2323 -1159
rect -2189 -1165 -2131 -1159
rect -1997 -1165 -1939 -1159
rect -1805 -1165 -1747 -1159
rect -1613 -1165 -1555 -1159
rect -1421 -1165 -1363 -1159
rect -1229 -1165 -1171 -1159
rect -1037 -1165 -979 -1159
rect -845 -1165 -787 -1159
rect -653 -1165 -595 -1159
rect -461 -1165 -403 -1159
rect -269 -1165 -211 -1159
rect -77 -1165 -19 -1159
rect 115 -1165 173 -1159
rect 307 -1165 365 -1159
rect 499 -1165 557 -1159
rect 691 -1165 749 -1159
rect 883 -1165 941 -1159
rect 1075 -1165 1133 -1159
rect 1267 -1165 1325 -1159
rect 1459 -1165 1517 -1159
rect 1651 -1165 1709 -1159
rect 1843 -1165 1901 -1159
rect 2035 -1165 2093 -1159
rect 2227 -1165 2285 -1159
rect -2381 -1199 -2369 -1165
rect -2189 -1199 -2177 -1165
rect -1997 -1199 -1985 -1165
rect -1805 -1199 -1793 -1165
rect -1613 -1199 -1601 -1165
rect -1421 -1199 -1409 -1165
rect -1229 -1199 -1217 -1165
rect -1037 -1199 -1025 -1165
rect -845 -1199 -833 -1165
rect -653 -1199 -641 -1165
rect -461 -1199 -449 -1165
rect -269 -1199 -257 -1165
rect -77 -1199 -65 -1165
rect 115 -1199 127 -1165
rect 307 -1199 319 -1165
rect 499 -1199 511 -1165
rect 691 -1199 703 -1165
rect 883 -1199 895 -1165
rect 1075 -1199 1087 -1165
rect 1267 -1199 1279 -1165
rect 1459 -1199 1471 -1165
rect 1651 -1199 1663 -1165
rect 1843 -1199 1855 -1165
rect 2035 -1199 2047 -1165
rect 2227 -1199 2239 -1165
rect -2381 -1205 -2323 -1199
rect -2189 -1205 -2131 -1199
rect -1997 -1205 -1939 -1199
rect -1805 -1205 -1747 -1199
rect -1613 -1205 -1555 -1199
rect -1421 -1205 -1363 -1199
rect -1229 -1205 -1171 -1199
rect -1037 -1205 -979 -1199
rect -845 -1205 -787 -1199
rect -653 -1205 -595 -1199
rect -461 -1205 -403 -1199
rect -269 -1205 -211 -1199
rect -77 -1205 -19 -1199
rect 115 -1205 173 -1199
rect 307 -1205 365 -1199
rect 499 -1205 557 -1199
rect 691 -1205 749 -1199
rect 883 -1205 941 -1199
rect 1075 -1205 1133 -1199
rect 1267 -1205 1325 -1199
rect 1459 -1205 1517 -1199
rect 1651 -1205 1709 -1199
rect 1843 -1205 1901 -1199
rect 2035 -1205 2093 -1199
rect 2227 -1205 2285 -1199
<< pwell >>
rect -2567 -1337 2567 1337
<< nmos >>
rect -2367 727 -2337 1127
rect -2271 727 -2241 1127
rect -2175 727 -2145 1127
rect -2079 727 -2049 1127
rect -1983 727 -1953 1127
rect -1887 727 -1857 1127
rect -1791 727 -1761 1127
rect -1695 727 -1665 1127
rect -1599 727 -1569 1127
rect -1503 727 -1473 1127
rect -1407 727 -1377 1127
rect -1311 727 -1281 1127
rect -1215 727 -1185 1127
rect -1119 727 -1089 1127
rect -1023 727 -993 1127
rect -927 727 -897 1127
rect -831 727 -801 1127
rect -735 727 -705 1127
rect -639 727 -609 1127
rect -543 727 -513 1127
rect -447 727 -417 1127
rect -351 727 -321 1127
rect -255 727 -225 1127
rect -159 727 -129 1127
rect -63 727 -33 1127
rect 33 727 63 1127
rect 129 727 159 1127
rect 225 727 255 1127
rect 321 727 351 1127
rect 417 727 447 1127
rect 513 727 543 1127
rect 609 727 639 1127
rect 705 727 735 1127
rect 801 727 831 1127
rect 897 727 927 1127
rect 993 727 1023 1127
rect 1089 727 1119 1127
rect 1185 727 1215 1127
rect 1281 727 1311 1127
rect 1377 727 1407 1127
rect 1473 727 1503 1127
rect 1569 727 1599 1127
rect 1665 727 1695 1127
rect 1761 727 1791 1127
rect 1857 727 1887 1127
rect 1953 727 1983 1127
rect 2049 727 2079 1127
rect 2145 727 2175 1127
rect 2241 727 2271 1127
rect 2337 727 2367 1127
rect -2367 109 -2337 509
rect -2271 109 -2241 509
rect -2175 109 -2145 509
rect -2079 109 -2049 509
rect -1983 109 -1953 509
rect -1887 109 -1857 509
rect -1791 109 -1761 509
rect -1695 109 -1665 509
rect -1599 109 -1569 509
rect -1503 109 -1473 509
rect -1407 109 -1377 509
rect -1311 109 -1281 509
rect -1215 109 -1185 509
rect -1119 109 -1089 509
rect -1023 109 -993 509
rect -927 109 -897 509
rect -831 109 -801 509
rect -735 109 -705 509
rect -639 109 -609 509
rect -543 109 -513 509
rect -447 109 -417 509
rect -351 109 -321 509
rect -255 109 -225 509
rect -159 109 -129 509
rect -63 109 -33 509
rect 33 109 63 509
rect 129 109 159 509
rect 225 109 255 509
rect 321 109 351 509
rect 417 109 447 509
rect 513 109 543 509
rect 609 109 639 509
rect 705 109 735 509
rect 801 109 831 509
rect 897 109 927 509
rect 993 109 1023 509
rect 1089 109 1119 509
rect 1185 109 1215 509
rect 1281 109 1311 509
rect 1377 109 1407 509
rect 1473 109 1503 509
rect 1569 109 1599 509
rect 1665 109 1695 509
rect 1761 109 1791 509
rect 1857 109 1887 509
rect 1953 109 1983 509
rect 2049 109 2079 509
rect 2145 109 2175 509
rect 2241 109 2271 509
rect 2337 109 2367 509
rect -2367 -509 -2337 -109
rect -2271 -509 -2241 -109
rect -2175 -509 -2145 -109
rect -2079 -509 -2049 -109
rect -1983 -509 -1953 -109
rect -1887 -509 -1857 -109
rect -1791 -509 -1761 -109
rect -1695 -509 -1665 -109
rect -1599 -509 -1569 -109
rect -1503 -509 -1473 -109
rect -1407 -509 -1377 -109
rect -1311 -509 -1281 -109
rect -1215 -509 -1185 -109
rect -1119 -509 -1089 -109
rect -1023 -509 -993 -109
rect -927 -509 -897 -109
rect -831 -509 -801 -109
rect -735 -509 -705 -109
rect -639 -509 -609 -109
rect -543 -509 -513 -109
rect -447 -509 -417 -109
rect -351 -509 -321 -109
rect -255 -509 -225 -109
rect -159 -509 -129 -109
rect -63 -509 -33 -109
rect 33 -509 63 -109
rect 129 -509 159 -109
rect 225 -509 255 -109
rect 321 -509 351 -109
rect 417 -509 447 -109
rect 513 -509 543 -109
rect 609 -509 639 -109
rect 705 -509 735 -109
rect 801 -509 831 -109
rect 897 -509 927 -109
rect 993 -509 1023 -109
rect 1089 -509 1119 -109
rect 1185 -509 1215 -109
rect 1281 -509 1311 -109
rect 1377 -509 1407 -109
rect 1473 -509 1503 -109
rect 1569 -509 1599 -109
rect 1665 -509 1695 -109
rect 1761 -509 1791 -109
rect 1857 -509 1887 -109
rect 1953 -509 1983 -109
rect 2049 -509 2079 -109
rect 2145 -509 2175 -109
rect 2241 -509 2271 -109
rect 2337 -509 2367 -109
rect -2367 -1127 -2337 -727
rect -2271 -1127 -2241 -727
rect -2175 -1127 -2145 -727
rect -2079 -1127 -2049 -727
rect -1983 -1127 -1953 -727
rect -1887 -1127 -1857 -727
rect -1791 -1127 -1761 -727
rect -1695 -1127 -1665 -727
rect -1599 -1127 -1569 -727
rect -1503 -1127 -1473 -727
rect -1407 -1127 -1377 -727
rect -1311 -1127 -1281 -727
rect -1215 -1127 -1185 -727
rect -1119 -1127 -1089 -727
rect -1023 -1127 -993 -727
rect -927 -1127 -897 -727
rect -831 -1127 -801 -727
rect -735 -1127 -705 -727
rect -639 -1127 -609 -727
rect -543 -1127 -513 -727
rect -447 -1127 -417 -727
rect -351 -1127 -321 -727
rect -255 -1127 -225 -727
rect -159 -1127 -129 -727
rect -63 -1127 -33 -727
rect 33 -1127 63 -727
rect 129 -1127 159 -727
rect 225 -1127 255 -727
rect 321 -1127 351 -727
rect 417 -1127 447 -727
rect 513 -1127 543 -727
rect 609 -1127 639 -727
rect 705 -1127 735 -727
rect 801 -1127 831 -727
rect 897 -1127 927 -727
rect 993 -1127 1023 -727
rect 1089 -1127 1119 -727
rect 1185 -1127 1215 -727
rect 1281 -1127 1311 -727
rect 1377 -1127 1407 -727
rect 1473 -1127 1503 -727
rect 1569 -1127 1599 -727
rect 1665 -1127 1695 -727
rect 1761 -1127 1791 -727
rect 1857 -1127 1887 -727
rect 1953 -1127 1983 -727
rect 2049 -1127 2079 -727
rect 2145 -1127 2175 -727
rect 2241 -1127 2271 -727
rect 2337 -1127 2367 -727
<< ndiff >>
rect -2429 1115 -2367 1127
rect -2429 739 -2417 1115
rect -2383 739 -2367 1115
rect -2429 727 -2367 739
rect -2337 1115 -2271 1127
rect -2337 739 -2321 1115
rect -2287 739 -2271 1115
rect -2337 727 -2271 739
rect -2241 1115 -2175 1127
rect -2241 739 -2225 1115
rect -2191 739 -2175 1115
rect -2241 727 -2175 739
rect -2145 1115 -2079 1127
rect -2145 739 -2129 1115
rect -2095 739 -2079 1115
rect -2145 727 -2079 739
rect -2049 1115 -1983 1127
rect -2049 739 -2033 1115
rect -1999 739 -1983 1115
rect -2049 727 -1983 739
rect -1953 1115 -1887 1127
rect -1953 739 -1937 1115
rect -1903 739 -1887 1115
rect -1953 727 -1887 739
rect -1857 1115 -1791 1127
rect -1857 739 -1841 1115
rect -1807 739 -1791 1115
rect -1857 727 -1791 739
rect -1761 1115 -1695 1127
rect -1761 739 -1745 1115
rect -1711 739 -1695 1115
rect -1761 727 -1695 739
rect -1665 1115 -1599 1127
rect -1665 739 -1649 1115
rect -1615 739 -1599 1115
rect -1665 727 -1599 739
rect -1569 1115 -1503 1127
rect -1569 739 -1553 1115
rect -1519 739 -1503 1115
rect -1569 727 -1503 739
rect -1473 1115 -1407 1127
rect -1473 739 -1457 1115
rect -1423 739 -1407 1115
rect -1473 727 -1407 739
rect -1377 1115 -1311 1127
rect -1377 739 -1361 1115
rect -1327 739 -1311 1115
rect -1377 727 -1311 739
rect -1281 1115 -1215 1127
rect -1281 739 -1265 1115
rect -1231 739 -1215 1115
rect -1281 727 -1215 739
rect -1185 1115 -1119 1127
rect -1185 739 -1169 1115
rect -1135 739 -1119 1115
rect -1185 727 -1119 739
rect -1089 1115 -1023 1127
rect -1089 739 -1073 1115
rect -1039 739 -1023 1115
rect -1089 727 -1023 739
rect -993 1115 -927 1127
rect -993 739 -977 1115
rect -943 739 -927 1115
rect -993 727 -927 739
rect -897 1115 -831 1127
rect -897 739 -881 1115
rect -847 739 -831 1115
rect -897 727 -831 739
rect -801 1115 -735 1127
rect -801 739 -785 1115
rect -751 739 -735 1115
rect -801 727 -735 739
rect -705 1115 -639 1127
rect -705 739 -689 1115
rect -655 739 -639 1115
rect -705 727 -639 739
rect -609 1115 -543 1127
rect -609 739 -593 1115
rect -559 739 -543 1115
rect -609 727 -543 739
rect -513 1115 -447 1127
rect -513 739 -497 1115
rect -463 739 -447 1115
rect -513 727 -447 739
rect -417 1115 -351 1127
rect -417 739 -401 1115
rect -367 739 -351 1115
rect -417 727 -351 739
rect -321 1115 -255 1127
rect -321 739 -305 1115
rect -271 739 -255 1115
rect -321 727 -255 739
rect -225 1115 -159 1127
rect -225 739 -209 1115
rect -175 739 -159 1115
rect -225 727 -159 739
rect -129 1115 -63 1127
rect -129 739 -113 1115
rect -79 739 -63 1115
rect -129 727 -63 739
rect -33 1115 33 1127
rect -33 739 -17 1115
rect 17 739 33 1115
rect -33 727 33 739
rect 63 1115 129 1127
rect 63 739 79 1115
rect 113 739 129 1115
rect 63 727 129 739
rect 159 1115 225 1127
rect 159 739 175 1115
rect 209 739 225 1115
rect 159 727 225 739
rect 255 1115 321 1127
rect 255 739 271 1115
rect 305 739 321 1115
rect 255 727 321 739
rect 351 1115 417 1127
rect 351 739 367 1115
rect 401 739 417 1115
rect 351 727 417 739
rect 447 1115 513 1127
rect 447 739 463 1115
rect 497 739 513 1115
rect 447 727 513 739
rect 543 1115 609 1127
rect 543 739 559 1115
rect 593 739 609 1115
rect 543 727 609 739
rect 639 1115 705 1127
rect 639 739 655 1115
rect 689 739 705 1115
rect 639 727 705 739
rect 735 1115 801 1127
rect 735 739 751 1115
rect 785 739 801 1115
rect 735 727 801 739
rect 831 1115 897 1127
rect 831 739 847 1115
rect 881 739 897 1115
rect 831 727 897 739
rect 927 1115 993 1127
rect 927 739 943 1115
rect 977 739 993 1115
rect 927 727 993 739
rect 1023 1115 1089 1127
rect 1023 739 1039 1115
rect 1073 739 1089 1115
rect 1023 727 1089 739
rect 1119 1115 1185 1127
rect 1119 739 1135 1115
rect 1169 739 1185 1115
rect 1119 727 1185 739
rect 1215 1115 1281 1127
rect 1215 739 1231 1115
rect 1265 739 1281 1115
rect 1215 727 1281 739
rect 1311 1115 1377 1127
rect 1311 739 1327 1115
rect 1361 739 1377 1115
rect 1311 727 1377 739
rect 1407 1115 1473 1127
rect 1407 739 1423 1115
rect 1457 739 1473 1115
rect 1407 727 1473 739
rect 1503 1115 1569 1127
rect 1503 739 1519 1115
rect 1553 739 1569 1115
rect 1503 727 1569 739
rect 1599 1115 1665 1127
rect 1599 739 1615 1115
rect 1649 739 1665 1115
rect 1599 727 1665 739
rect 1695 1115 1761 1127
rect 1695 739 1711 1115
rect 1745 739 1761 1115
rect 1695 727 1761 739
rect 1791 1115 1857 1127
rect 1791 739 1807 1115
rect 1841 739 1857 1115
rect 1791 727 1857 739
rect 1887 1115 1953 1127
rect 1887 739 1903 1115
rect 1937 739 1953 1115
rect 1887 727 1953 739
rect 1983 1115 2049 1127
rect 1983 739 1999 1115
rect 2033 739 2049 1115
rect 1983 727 2049 739
rect 2079 1115 2145 1127
rect 2079 739 2095 1115
rect 2129 739 2145 1115
rect 2079 727 2145 739
rect 2175 1115 2241 1127
rect 2175 739 2191 1115
rect 2225 739 2241 1115
rect 2175 727 2241 739
rect 2271 1115 2337 1127
rect 2271 739 2287 1115
rect 2321 739 2337 1115
rect 2271 727 2337 739
rect 2367 1115 2429 1127
rect 2367 739 2383 1115
rect 2417 739 2429 1115
rect 2367 727 2429 739
rect -2429 497 -2367 509
rect -2429 121 -2417 497
rect -2383 121 -2367 497
rect -2429 109 -2367 121
rect -2337 497 -2271 509
rect -2337 121 -2321 497
rect -2287 121 -2271 497
rect -2337 109 -2271 121
rect -2241 497 -2175 509
rect -2241 121 -2225 497
rect -2191 121 -2175 497
rect -2241 109 -2175 121
rect -2145 497 -2079 509
rect -2145 121 -2129 497
rect -2095 121 -2079 497
rect -2145 109 -2079 121
rect -2049 497 -1983 509
rect -2049 121 -2033 497
rect -1999 121 -1983 497
rect -2049 109 -1983 121
rect -1953 497 -1887 509
rect -1953 121 -1937 497
rect -1903 121 -1887 497
rect -1953 109 -1887 121
rect -1857 497 -1791 509
rect -1857 121 -1841 497
rect -1807 121 -1791 497
rect -1857 109 -1791 121
rect -1761 497 -1695 509
rect -1761 121 -1745 497
rect -1711 121 -1695 497
rect -1761 109 -1695 121
rect -1665 497 -1599 509
rect -1665 121 -1649 497
rect -1615 121 -1599 497
rect -1665 109 -1599 121
rect -1569 497 -1503 509
rect -1569 121 -1553 497
rect -1519 121 -1503 497
rect -1569 109 -1503 121
rect -1473 497 -1407 509
rect -1473 121 -1457 497
rect -1423 121 -1407 497
rect -1473 109 -1407 121
rect -1377 497 -1311 509
rect -1377 121 -1361 497
rect -1327 121 -1311 497
rect -1377 109 -1311 121
rect -1281 497 -1215 509
rect -1281 121 -1265 497
rect -1231 121 -1215 497
rect -1281 109 -1215 121
rect -1185 497 -1119 509
rect -1185 121 -1169 497
rect -1135 121 -1119 497
rect -1185 109 -1119 121
rect -1089 497 -1023 509
rect -1089 121 -1073 497
rect -1039 121 -1023 497
rect -1089 109 -1023 121
rect -993 497 -927 509
rect -993 121 -977 497
rect -943 121 -927 497
rect -993 109 -927 121
rect -897 497 -831 509
rect -897 121 -881 497
rect -847 121 -831 497
rect -897 109 -831 121
rect -801 497 -735 509
rect -801 121 -785 497
rect -751 121 -735 497
rect -801 109 -735 121
rect -705 497 -639 509
rect -705 121 -689 497
rect -655 121 -639 497
rect -705 109 -639 121
rect -609 497 -543 509
rect -609 121 -593 497
rect -559 121 -543 497
rect -609 109 -543 121
rect -513 497 -447 509
rect -513 121 -497 497
rect -463 121 -447 497
rect -513 109 -447 121
rect -417 497 -351 509
rect -417 121 -401 497
rect -367 121 -351 497
rect -417 109 -351 121
rect -321 497 -255 509
rect -321 121 -305 497
rect -271 121 -255 497
rect -321 109 -255 121
rect -225 497 -159 509
rect -225 121 -209 497
rect -175 121 -159 497
rect -225 109 -159 121
rect -129 497 -63 509
rect -129 121 -113 497
rect -79 121 -63 497
rect -129 109 -63 121
rect -33 497 33 509
rect -33 121 -17 497
rect 17 121 33 497
rect -33 109 33 121
rect 63 497 129 509
rect 63 121 79 497
rect 113 121 129 497
rect 63 109 129 121
rect 159 497 225 509
rect 159 121 175 497
rect 209 121 225 497
rect 159 109 225 121
rect 255 497 321 509
rect 255 121 271 497
rect 305 121 321 497
rect 255 109 321 121
rect 351 497 417 509
rect 351 121 367 497
rect 401 121 417 497
rect 351 109 417 121
rect 447 497 513 509
rect 447 121 463 497
rect 497 121 513 497
rect 447 109 513 121
rect 543 497 609 509
rect 543 121 559 497
rect 593 121 609 497
rect 543 109 609 121
rect 639 497 705 509
rect 639 121 655 497
rect 689 121 705 497
rect 639 109 705 121
rect 735 497 801 509
rect 735 121 751 497
rect 785 121 801 497
rect 735 109 801 121
rect 831 497 897 509
rect 831 121 847 497
rect 881 121 897 497
rect 831 109 897 121
rect 927 497 993 509
rect 927 121 943 497
rect 977 121 993 497
rect 927 109 993 121
rect 1023 497 1089 509
rect 1023 121 1039 497
rect 1073 121 1089 497
rect 1023 109 1089 121
rect 1119 497 1185 509
rect 1119 121 1135 497
rect 1169 121 1185 497
rect 1119 109 1185 121
rect 1215 497 1281 509
rect 1215 121 1231 497
rect 1265 121 1281 497
rect 1215 109 1281 121
rect 1311 497 1377 509
rect 1311 121 1327 497
rect 1361 121 1377 497
rect 1311 109 1377 121
rect 1407 497 1473 509
rect 1407 121 1423 497
rect 1457 121 1473 497
rect 1407 109 1473 121
rect 1503 497 1569 509
rect 1503 121 1519 497
rect 1553 121 1569 497
rect 1503 109 1569 121
rect 1599 497 1665 509
rect 1599 121 1615 497
rect 1649 121 1665 497
rect 1599 109 1665 121
rect 1695 497 1761 509
rect 1695 121 1711 497
rect 1745 121 1761 497
rect 1695 109 1761 121
rect 1791 497 1857 509
rect 1791 121 1807 497
rect 1841 121 1857 497
rect 1791 109 1857 121
rect 1887 497 1953 509
rect 1887 121 1903 497
rect 1937 121 1953 497
rect 1887 109 1953 121
rect 1983 497 2049 509
rect 1983 121 1999 497
rect 2033 121 2049 497
rect 1983 109 2049 121
rect 2079 497 2145 509
rect 2079 121 2095 497
rect 2129 121 2145 497
rect 2079 109 2145 121
rect 2175 497 2241 509
rect 2175 121 2191 497
rect 2225 121 2241 497
rect 2175 109 2241 121
rect 2271 497 2337 509
rect 2271 121 2287 497
rect 2321 121 2337 497
rect 2271 109 2337 121
rect 2367 497 2429 509
rect 2367 121 2383 497
rect 2417 121 2429 497
rect 2367 109 2429 121
rect -2429 -121 -2367 -109
rect -2429 -497 -2417 -121
rect -2383 -497 -2367 -121
rect -2429 -509 -2367 -497
rect -2337 -121 -2271 -109
rect -2337 -497 -2321 -121
rect -2287 -497 -2271 -121
rect -2337 -509 -2271 -497
rect -2241 -121 -2175 -109
rect -2241 -497 -2225 -121
rect -2191 -497 -2175 -121
rect -2241 -509 -2175 -497
rect -2145 -121 -2079 -109
rect -2145 -497 -2129 -121
rect -2095 -497 -2079 -121
rect -2145 -509 -2079 -497
rect -2049 -121 -1983 -109
rect -2049 -497 -2033 -121
rect -1999 -497 -1983 -121
rect -2049 -509 -1983 -497
rect -1953 -121 -1887 -109
rect -1953 -497 -1937 -121
rect -1903 -497 -1887 -121
rect -1953 -509 -1887 -497
rect -1857 -121 -1791 -109
rect -1857 -497 -1841 -121
rect -1807 -497 -1791 -121
rect -1857 -509 -1791 -497
rect -1761 -121 -1695 -109
rect -1761 -497 -1745 -121
rect -1711 -497 -1695 -121
rect -1761 -509 -1695 -497
rect -1665 -121 -1599 -109
rect -1665 -497 -1649 -121
rect -1615 -497 -1599 -121
rect -1665 -509 -1599 -497
rect -1569 -121 -1503 -109
rect -1569 -497 -1553 -121
rect -1519 -497 -1503 -121
rect -1569 -509 -1503 -497
rect -1473 -121 -1407 -109
rect -1473 -497 -1457 -121
rect -1423 -497 -1407 -121
rect -1473 -509 -1407 -497
rect -1377 -121 -1311 -109
rect -1377 -497 -1361 -121
rect -1327 -497 -1311 -121
rect -1377 -509 -1311 -497
rect -1281 -121 -1215 -109
rect -1281 -497 -1265 -121
rect -1231 -497 -1215 -121
rect -1281 -509 -1215 -497
rect -1185 -121 -1119 -109
rect -1185 -497 -1169 -121
rect -1135 -497 -1119 -121
rect -1185 -509 -1119 -497
rect -1089 -121 -1023 -109
rect -1089 -497 -1073 -121
rect -1039 -497 -1023 -121
rect -1089 -509 -1023 -497
rect -993 -121 -927 -109
rect -993 -497 -977 -121
rect -943 -497 -927 -121
rect -993 -509 -927 -497
rect -897 -121 -831 -109
rect -897 -497 -881 -121
rect -847 -497 -831 -121
rect -897 -509 -831 -497
rect -801 -121 -735 -109
rect -801 -497 -785 -121
rect -751 -497 -735 -121
rect -801 -509 -735 -497
rect -705 -121 -639 -109
rect -705 -497 -689 -121
rect -655 -497 -639 -121
rect -705 -509 -639 -497
rect -609 -121 -543 -109
rect -609 -497 -593 -121
rect -559 -497 -543 -121
rect -609 -509 -543 -497
rect -513 -121 -447 -109
rect -513 -497 -497 -121
rect -463 -497 -447 -121
rect -513 -509 -447 -497
rect -417 -121 -351 -109
rect -417 -497 -401 -121
rect -367 -497 -351 -121
rect -417 -509 -351 -497
rect -321 -121 -255 -109
rect -321 -497 -305 -121
rect -271 -497 -255 -121
rect -321 -509 -255 -497
rect -225 -121 -159 -109
rect -225 -497 -209 -121
rect -175 -497 -159 -121
rect -225 -509 -159 -497
rect -129 -121 -63 -109
rect -129 -497 -113 -121
rect -79 -497 -63 -121
rect -129 -509 -63 -497
rect -33 -121 33 -109
rect -33 -497 -17 -121
rect 17 -497 33 -121
rect -33 -509 33 -497
rect 63 -121 129 -109
rect 63 -497 79 -121
rect 113 -497 129 -121
rect 63 -509 129 -497
rect 159 -121 225 -109
rect 159 -497 175 -121
rect 209 -497 225 -121
rect 159 -509 225 -497
rect 255 -121 321 -109
rect 255 -497 271 -121
rect 305 -497 321 -121
rect 255 -509 321 -497
rect 351 -121 417 -109
rect 351 -497 367 -121
rect 401 -497 417 -121
rect 351 -509 417 -497
rect 447 -121 513 -109
rect 447 -497 463 -121
rect 497 -497 513 -121
rect 447 -509 513 -497
rect 543 -121 609 -109
rect 543 -497 559 -121
rect 593 -497 609 -121
rect 543 -509 609 -497
rect 639 -121 705 -109
rect 639 -497 655 -121
rect 689 -497 705 -121
rect 639 -509 705 -497
rect 735 -121 801 -109
rect 735 -497 751 -121
rect 785 -497 801 -121
rect 735 -509 801 -497
rect 831 -121 897 -109
rect 831 -497 847 -121
rect 881 -497 897 -121
rect 831 -509 897 -497
rect 927 -121 993 -109
rect 927 -497 943 -121
rect 977 -497 993 -121
rect 927 -509 993 -497
rect 1023 -121 1089 -109
rect 1023 -497 1039 -121
rect 1073 -497 1089 -121
rect 1023 -509 1089 -497
rect 1119 -121 1185 -109
rect 1119 -497 1135 -121
rect 1169 -497 1185 -121
rect 1119 -509 1185 -497
rect 1215 -121 1281 -109
rect 1215 -497 1231 -121
rect 1265 -497 1281 -121
rect 1215 -509 1281 -497
rect 1311 -121 1377 -109
rect 1311 -497 1327 -121
rect 1361 -497 1377 -121
rect 1311 -509 1377 -497
rect 1407 -121 1473 -109
rect 1407 -497 1423 -121
rect 1457 -497 1473 -121
rect 1407 -509 1473 -497
rect 1503 -121 1569 -109
rect 1503 -497 1519 -121
rect 1553 -497 1569 -121
rect 1503 -509 1569 -497
rect 1599 -121 1665 -109
rect 1599 -497 1615 -121
rect 1649 -497 1665 -121
rect 1599 -509 1665 -497
rect 1695 -121 1761 -109
rect 1695 -497 1711 -121
rect 1745 -497 1761 -121
rect 1695 -509 1761 -497
rect 1791 -121 1857 -109
rect 1791 -497 1807 -121
rect 1841 -497 1857 -121
rect 1791 -509 1857 -497
rect 1887 -121 1953 -109
rect 1887 -497 1903 -121
rect 1937 -497 1953 -121
rect 1887 -509 1953 -497
rect 1983 -121 2049 -109
rect 1983 -497 1999 -121
rect 2033 -497 2049 -121
rect 1983 -509 2049 -497
rect 2079 -121 2145 -109
rect 2079 -497 2095 -121
rect 2129 -497 2145 -121
rect 2079 -509 2145 -497
rect 2175 -121 2241 -109
rect 2175 -497 2191 -121
rect 2225 -497 2241 -121
rect 2175 -509 2241 -497
rect 2271 -121 2337 -109
rect 2271 -497 2287 -121
rect 2321 -497 2337 -121
rect 2271 -509 2337 -497
rect 2367 -121 2429 -109
rect 2367 -497 2383 -121
rect 2417 -497 2429 -121
rect 2367 -509 2429 -497
rect -2429 -739 -2367 -727
rect -2429 -1115 -2417 -739
rect -2383 -1115 -2367 -739
rect -2429 -1127 -2367 -1115
rect -2337 -739 -2271 -727
rect -2337 -1115 -2321 -739
rect -2287 -1115 -2271 -739
rect -2337 -1127 -2271 -1115
rect -2241 -739 -2175 -727
rect -2241 -1115 -2225 -739
rect -2191 -1115 -2175 -739
rect -2241 -1127 -2175 -1115
rect -2145 -739 -2079 -727
rect -2145 -1115 -2129 -739
rect -2095 -1115 -2079 -739
rect -2145 -1127 -2079 -1115
rect -2049 -739 -1983 -727
rect -2049 -1115 -2033 -739
rect -1999 -1115 -1983 -739
rect -2049 -1127 -1983 -1115
rect -1953 -739 -1887 -727
rect -1953 -1115 -1937 -739
rect -1903 -1115 -1887 -739
rect -1953 -1127 -1887 -1115
rect -1857 -739 -1791 -727
rect -1857 -1115 -1841 -739
rect -1807 -1115 -1791 -739
rect -1857 -1127 -1791 -1115
rect -1761 -739 -1695 -727
rect -1761 -1115 -1745 -739
rect -1711 -1115 -1695 -739
rect -1761 -1127 -1695 -1115
rect -1665 -739 -1599 -727
rect -1665 -1115 -1649 -739
rect -1615 -1115 -1599 -739
rect -1665 -1127 -1599 -1115
rect -1569 -739 -1503 -727
rect -1569 -1115 -1553 -739
rect -1519 -1115 -1503 -739
rect -1569 -1127 -1503 -1115
rect -1473 -739 -1407 -727
rect -1473 -1115 -1457 -739
rect -1423 -1115 -1407 -739
rect -1473 -1127 -1407 -1115
rect -1377 -739 -1311 -727
rect -1377 -1115 -1361 -739
rect -1327 -1115 -1311 -739
rect -1377 -1127 -1311 -1115
rect -1281 -739 -1215 -727
rect -1281 -1115 -1265 -739
rect -1231 -1115 -1215 -739
rect -1281 -1127 -1215 -1115
rect -1185 -739 -1119 -727
rect -1185 -1115 -1169 -739
rect -1135 -1115 -1119 -739
rect -1185 -1127 -1119 -1115
rect -1089 -739 -1023 -727
rect -1089 -1115 -1073 -739
rect -1039 -1115 -1023 -739
rect -1089 -1127 -1023 -1115
rect -993 -739 -927 -727
rect -993 -1115 -977 -739
rect -943 -1115 -927 -739
rect -993 -1127 -927 -1115
rect -897 -739 -831 -727
rect -897 -1115 -881 -739
rect -847 -1115 -831 -739
rect -897 -1127 -831 -1115
rect -801 -739 -735 -727
rect -801 -1115 -785 -739
rect -751 -1115 -735 -739
rect -801 -1127 -735 -1115
rect -705 -739 -639 -727
rect -705 -1115 -689 -739
rect -655 -1115 -639 -739
rect -705 -1127 -639 -1115
rect -609 -739 -543 -727
rect -609 -1115 -593 -739
rect -559 -1115 -543 -739
rect -609 -1127 -543 -1115
rect -513 -739 -447 -727
rect -513 -1115 -497 -739
rect -463 -1115 -447 -739
rect -513 -1127 -447 -1115
rect -417 -739 -351 -727
rect -417 -1115 -401 -739
rect -367 -1115 -351 -739
rect -417 -1127 -351 -1115
rect -321 -739 -255 -727
rect -321 -1115 -305 -739
rect -271 -1115 -255 -739
rect -321 -1127 -255 -1115
rect -225 -739 -159 -727
rect -225 -1115 -209 -739
rect -175 -1115 -159 -739
rect -225 -1127 -159 -1115
rect -129 -739 -63 -727
rect -129 -1115 -113 -739
rect -79 -1115 -63 -739
rect -129 -1127 -63 -1115
rect -33 -739 33 -727
rect -33 -1115 -17 -739
rect 17 -1115 33 -739
rect -33 -1127 33 -1115
rect 63 -739 129 -727
rect 63 -1115 79 -739
rect 113 -1115 129 -739
rect 63 -1127 129 -1115
rect 159 -739 225 -727
rect 159 -1115 175 -739
rect 209 -1115 225 -739
rect 159 -1127 225 -1115
rect 255 -739 321 -727
rect 255 -1115 271 -739
rect 305 -1115 321 -739
rect 255 -1127 321 -1115
rect 351 -739 417 -727
rect 351 -1115 367 -739
rect 401 -1115 417 -739
rect 351 -1127 417 -1115
rect 447 -739 513 -727
rect 447 -1115 463 -739
rect 497 -1115 513 -739
rect 447 -1127 513 -1115
rect 543 -739 609 -727
rect 543 -1115 559 -739
rect 593 -1115 609 -739
rect 543 -1127 609 -1115
rect 639 -739 705 -727
rect 639 -1115 655 -739
rect 689 -1115 705 -739
rect 639 -1127 705 -1115
rect 735 -739 801 -727
rect 735 -1115 751 -739
rect 785 -1115 801 -739
rect 735 -1127 801 -1115
rect 831 -739 897 -727
rect 831 -1115 847 -739
rect 881 -1115 897 -739
rect 831 -1127 897 -1115
rect 927 -739 993 -727
rect 927 -1115 943 -739
rect 977 -1115 993 -739
rect 927 -1127 993 -1115
rect 1023 -739 1089 -727
rect 1023 -1115 1039 -739
rect 1073 -1115 1089 -739
rect 1023 -1127 1089 -1115
rect 1119 -739 1185 -727
rect 1119 -1115 1135 -739
rect 1169 -1115 1185 -739
rect 1119 -1127 1185 -1115
rect 1215 -739 1281 -727
rect 1215 -1115 1231 -739
rect 1265 -1115 1281 -739
rect 1215 -1127 1281 -1115
rect 1311 -739 1377 -727
rect 1311 -1115 1327 -739
rect 1361 -1115 1377 -739
rect 1311 -1127 1377 -1115
rect 1407 -739 1473 -727
rect 1407 -1115 1423 -739
rect 1457 -1115 1473 -739
rect 1407 -1127 1473 -1115
rect 1503 -739 1569 -727
rect 1503 -1115 1519 -739
rect 1553 -1115 1569 -739
rect 1503 -1127 1569 -1115
rect 1599 -739 1665 -727
rect 1599 -1115 1615 -739
rect 1649 -1115 1665 -739
rect 1599 -1127 1665 -1115
rect 1695 -739 1761 -727
rect 1695 -1115 1711 -739
rect 1745 -1115 1761 -739
rect 1695 -1127 1761 -1115
rect 1791 -739 1857 -727
rect 1791 -1115 1807 -739
rect 1841 -1115 1857 -739
rect 1791 -1127 1857 -1115
rect 1887 -739 1953 -727
rect 1887 -1115 1903 -739
rect 1937 -1115 1953 -739
rect 1887 -1127 1953 -1115
rect 1983 -739 2049 -727
rect 1983 -1115 1999 -739
rect 2033 -1115 2049 -739
rect 1983 -1127 2049 -1115
rect 2079 -739 2145 -727
rect 2079 -1115 2095 -739
rect 2129 -1115 2145 -739
rect 2079 -1127 2145 -1115
rect 2175 -739 2241 -727
rect 2175 -1115 2191 -739
rect 2225 -1115 2241 -739
rect 2175 -1127 2241 -1115
rect 2271 -739 2337 -727
rect 2271 -1115 2287 -739
rect 2321 -1115 2337 -739
rect 2271 -1127 2337 -1115
rect 2367 -739 2429 -727
rect 2367 -1115 2383 -739
rect 2417 -1115 2429 -739
rect 2367 -1127 2429 -1115
<< ndiffc >>
rect -2417 739 -2383 1115
rect -2321 739 -2287 1115
rect -2225 739 -2191 1115
rect -2129 739 -2095 1115
rect -2033 739 -1999 1115
rect -1937 739 -1903 1115
rect -1841 739 -1807 1115
rect -1745 739 -1711 1115
rect -1649 739 -1615 1115
rect -1553 739 -1519 1115
rect -1457 739 -1423 1115
rect -1361 739 -1327 1115
rect -1265 739 -1231 1115
rect -1169 739 -1135 1115
rect -1073 739 -1039 1115
rect -977 739 -943 1115
rect -881 739 -847 1115
rect -785 739 -751 1115
rect -689 739 -655 1115
rect -593 739 -559 1115
rect -497 739 -463 1115
rect -401 739 -367 1115
rect -305 739 -271 1115
rect -209 739 -175 1115
rect -113 739 -79 1115
rect -17 739 17 1115
rect 79 739 113 1115
rect 175 739 209 1115
rect 271 739 305 1115
rect 367 739 401 1115
rect 463 739 497 1115
rect 559 739 593 1115
rect 655 739 689 1115
rect 751 739 785 1115
rect 847 739 881 1115
rect 943 739 977 1115
rect 1039 739 1073 1115
rect 1135 739 1169 1115
rect 1231 739 1265 1115
rect 1327 739 1361 1115
rect 1423 739 1457 1115
rect 1519 739 1553 1115
rect 1615 739 1649 1115
rect 1711 739 1745 1115
rect 1807 739 1841 1115
rect 1903 739 1937 1115
rect 1999 739 2033 1115
rect 2095 739 2129 1115
rect 2191 739 2225 1115
rect 2287 739 2321 1115
rect 2383 739 2417 1115
rect -2417 121 -2383 497
rect -2321 121 -2287 497
rect -2225 121 -2191 497
rect -2129 121 -2095 497
rect -2033 121 -1999 497
rect -1937 121 -1903 497
rect -1841 121 -1807 497
rect -1745 121 -1711 497
rect -1649 121 -1615 497
rect -1553 121 -1519 497
rect -1457 121 -1423 497
rect -1361 121 -1327 497
rect -1265 121 -1231 497
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect 1231 121 1265 497
rect 1327 121 1361 497
rect 1423 121 1457 497
rect 1519 121 1553 497
rect 1615 121 1649 497
rect 1711 121 1745 497
rect 1807 121 1841 497
rect 1903 121 1937 497
rect 1999 121 2033 497
rect 2095 121 2129 497
rect 2191 121 2225 497
rect 2287 121 2321 497
rect 2383 121 2417 497
rect -2417 -497 -2383 -121
rect -2321 -497 -2287 -121
rect -2225 -497 -2191 -121
rect -2129 -497 -2095 -121
rect -2033 -497 -1999 -121
rect -1937 -497 -1903 -121
rect -1841 -497 -1807 -121
rect -1745 -497 -1711 -121
rect -1649 -497 -1615 -121
rect -1553 -497 -1519 -121
rect -1457 -497 -1423 -121
rect -1361 -497 -1327 -121
rect -1265 -497 -1231 -121
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect 1231 -497 1265 -121
rect 1327 -497 1361 -121
rect 1423 -497 1457 -121
rect 1519 -497 1553 -121
rect 1615 -497 1649 -121
rect 1711 -497 1745 -121
rect 1807 -497 1841 -121
rect 1903 -497 1937 -121
rect 1999 -497 2033 -121
rect 2095 -497 2129 -121
rect 2191 -497 2225 -121
rect 2287 -497 2321 -121
rect 2383 -497 2417 -121
rect -2417 -1115 -2383 -739
rect -2321 -1115 -2287 -739
rect -2225 -1115 -2191 -739
rect -2129 -1115 -2095 -739
rect -2033 -1115 -1999 -739
rect -1937 -1115 -1903 -739
rect -1841 -1115 -1807 -739
rect -1745 -1115 -1711 -739
rect -1649 -1115 -1615 -739
rect -1553 -1115 -1519 -739
rect -1457 -1115 -1423 -739
rect -1361 -1115 -1327 -739
rect -1265 -1115 -1231 -739
rect -1169 -1115 -1135 -739
rect -1073 -1115 -1039 -739
rect -977 -1115 -943 -739
rect -881 -1115 -847 -739
rect -785 -1115 -751 -739
rect -689 -1115 -655 -739
rect -593 -1115 -559 -739
rect -497 -1115 -463 -739
rect -401 -1115 -367 -739
rect -305 -1115 -271 -739
rect -209 -1115 -175 -739
rect -113 -1115 -79 -739
rect -17 -1115 17 -739
rect 79 -1115 113 -739
rect 175 -1115 209 -739
rect 271 -1115 305 -739
rect 367 -1115 401 -739
rect 463 -1115 497 -739
rect 559 -1115 593 -739
rect 655 -1115 689 -739
rect 751 -1115 785 -739
rect 847 -1115 881 -739
rect 943 -1115 977 -739
rect 1039 -1115 1073 -739
rect 1135 -1115 1169 -739
rect 1231 -1115 1265 -739
rect 1327 -1115 1361 -739
rect 1423 -1115 1457 -739
rect 1519 -1115 1553 -739
rect 1615 -1115 1649 -739
rect 1711 -1115 1745 -739
rect 1807 -1115 1841 -739
rect 1903 -1115 1937 -739
rect 1999 -1115 2033 -739
rect 2095 -1115 2129 -739
rect 2191 -1115 2225 -739
rect 2287 -1115 2321 -739
rect 2383 -1115 2417 -739
<< psubdiff >>
rect -2531 1267 -2435 1301
rect 2435 1267 2531 1301
rect -2531 1205 -2497 1267
rect 2497 1205 2531 1267
rect -2531 -1267 -2497 -1205
rect 2497 -1267 2531 -1205
rect -2531 -1301 -2435 -1267
rect 2435 -1301 2531 -1267
<< psubdiffcont >>
rect -2435 1267 2435 1301
rect -2531 -1205 -2497 1205
rect 2497 -1205 2531 1205
rect -2435 -1301 2435 -1267
<< poly >>
rect -2385 1199 -2319 1215
rect -2385 1165 -2369 1199
rect -2335 1165 -2319 1199
rect -2385 1149 -2319 1165
rect -2193 1199 -2127 1215
rect -2193 1165 -2177 1199
rect -2143 1165 -2127 1199
rect -2367 1127 -2337 1149
rect -2271 1127 -2241 1153
rect -2193 1149 -2127 1165
rect -2001 1199 -1935 1215
rect -2001 1165 -1985 1199
rect -1951 1165 -1935 1199
rect -2175 1127 -2145 1149
rect -2079 1127 -2049 1153
rect -2001 1149 -1935 1165
rect -1809 1199 -1743 1215
rect -1809 1165 -1793 1199
rect -1759 1165 -1743 1199
rect -1983 1127 -1953 1149
rect -1887 1127 -1857 1153
rect -1809 1149 -1743 1165
rect -1617 1199 -1551 1215
rect -1617 1165 -1601 1199
rect -1567 1165 -1551 1199
rect -1791 1127 -1761 1149
rect -1695 1127 -1665 1153
rect -1617 1149 -1551 1165
rect -1425 1199 -1359 1215
rect -1425 1165 -1409 1199
rect -1375 1165 -1359 1199
rect -1599 1127 -1569 1149
rect -1503 1127 -1473 1153
rect -1425 1149 -1359 1165
rect -1233 1199 -1167 1215
rect -1233 1165 -1217 1199
rect -1183 1165 -1167 1199
rect -1407 1127 -1377 1149
rect -1311 1127 -1281 1153
rect -1233 1149 -1167 1165
rect -1041 1199 -975 1215
rect -1041 1165 -1025 1199
rect -991 1165 -975 1199
rect -1215 1127 -1185 1149
rect -1119 1127 -1089 1153
rect -1041 1149 -975 1165
rect -849 1199 -783 1215
rect -849 1165 -833 1199
rect -799 1165 -783 1199
rect -1023 1127 -993 1149
rect -927 1127 -897 1153
rect -849 1149 -783 1165
rect -657 1199 -591 1215
rect -657 1165 -641 1199
rect -607 1165 -591 1199
rect -831 1127 -801 1149
rect -735 1127 -705 1153
rect -657 1149 -591 1165
rect -465 1199 -399 1215
rect -465 1165 -449 1199
rect -415 1165 -399 1199
rect -639 1127 -609 1149
rect -543 1127 -513 1153
rect -465 1149 -399 1165
rect -273 1199 -207 1215
rect -273 1165 -257 1199
rect -223 1165 -207 1199
rect -447 1127 -417 1149
rect -351 1127 -321 1153
rect -273 1149 -207 1165
rect -81 1199 -15 1215
rect -81 1165 -65 1199
rect -31 1165 -15 1199
rect -255 1127 -225 1149
rect -159 1127 -129 1153
rect -81 1149 -15 1165
rect 111 1199 177 1215
rect 111 1165 127 1199
rect 161 1165 177 1199
rect -63 1127 -33 1149
rect 33 1127 63 1153
rect 111 1149 177 1165
rect 303 1199 369 1215
rect 303 1165 319 1199
rect 353 1165 369 1199
rect 129 1127 159 1149
rect 225 1127 255 1153
rect 303 1149 369 1165
rect 495 1199 561 1215
rect 495 1165 511 1199
rect 545 1165 561 1199
rect 321 1127 351 1149
rect 417 1127 447 1153
rect 495 1149 561 1165
rect 687 1199 753 1215
rect 687 1165 703 1199
rect 737 1165 753 1199
rect 513 1127 543 1149
rect 609 1127 639 1153
rect 687 1149 753 1165
rect 879 1199 945 1215
rect 879 1165 895 1199
rect 929 1165 945 1199
rect 705 1127 735 1149
rect 801 1127 831 1153
rect 879 1149 945 1165
rect 1071 1199 1137 1215
rect 1071 1165 1087 1199
rect 1121 1165 1137 1199
rect 897 1127 927 1149
rect 993 1127 1023 1153
rect 1071 1149 1137 1165
rect 1263 1199 1329 1215
rect 1263 1165 1279 1199
rect 1313 1165 1329 1199
rect 1089 1127 1119 1149
rect 1185 1127 1215 1153
rect 1263 1149 1329 1165
rect 1455 1199 1521 1215
rect 1455 1165 1471 1199
rect 1505 1165 1521 1199
rect 1281 1127 1311 1149
rect 1377 1127 1407 1153
rect 1455 1149 1521 1165
rect 1647 1199 1713 1215
rect 1647 1165 1663 1199
rect 1697 1165 1713 1199
rect 1473 1127 1503 1149
rect 1569 1127 1599 1153
rect 1647 1149 1713 1165
rect 1839 1199 1905 1215
rect 1839 1165 1855 1199
rect 1889 1165 1905 1199
rect 1665 1127 1695 1149
rect 1761 1127 1791 1153
rect 1839 1149 1905 1165
rect 2031 1199 2097 1215
rect 2031 1165 2047 1199
rect 2081 1165 2097 1199
rect 1857 1127 1887 1149
rect 1953 1127 1983 1153
rect 2031 1149 2097 1165
rect 2223 1199 2289 1215
rect 2223 1165 2239 1199
rect 2273 1165 2289 1199
rect 2049 1127 2079 1149
rect 2145 1127 2175 1153
rect 2223 1149 2289 1165
rect 2241 1127 2271 1149
rect 2337 1127 2367 1153
rect -2367 701 -2337 727
rect -2271 705 -2241 727
rect -2289 689 -2223 705
rect -2175 701 -2145 727
rect -2079 705 -2049 727
rect -2289 655 -2273 689
rect -2239 655 -2223 689
rect -2289 639 -2223 655
rect -2097 689 -2031 705
rect -1983 701 -1953 727
rect -1887 705 -1857 727
rect -2097 655 -2081 689
rect -2047 655 -2031 689
rect -2097 639 -2031 655
rect -1905 689 -1839 705
rect -1791 701 -1761 727
rect -1695 705 -1665 727
rect -1905 655 -1889 689
rect -1855 655 -1839 689
rect -1905 639 -1839 655
rect -1713 689 -1647 705
rect -1599 701 -1569 727
rect -1503 705 -1473 727
rect -1713 655 -1697 689
rect -1663 655 -1647 689
rect -1713 639 -1647 655
rect -1521 689 -1455 705
rect -1407 701 -1377 727
rect -1311 705 -1281 727
rect -1521 655 -1505 689
rect -1471 655 -1455 689
rect -1521 639 -1455 655
rect -1329 689 -1263 705
rect -1215 701 -1185 727
rect -1119 705 -1089 727
rect -1329 655 -1313 689
rect -1279 655 -1263 689
rect -1329 639 -1263 655
rect -1137 689 -1071 705
rect -1023 701 -993 727
rect -927 705 -897 727
rect -1137 655 -1121 689
rect -1087 655 -1071 689
rect -1137 639 -1071 655
rect -945 689 -879 705
rect -831 701 -801 727
rect -735 705 -705 727
rect -945 655 -929 689
rect -895 655 -879 689
rect -945 639 -879 655
rect -753 689 -687 705
rect -639 701 -609 727
rect -543 705 -513 727
rect -753 655 -737 689
rect -703 655 -687 689
rect -753 639 -687 655
rect -561 689 -495 705
rect -447 701 -417 727
rect -351 705 -321 727
rect -561 655 -545 689
rect -511 655 -495 689
rect -561 639 -495 655
rect -369 689 -303 705
rect -255 701 -225 727
rect -159 705 -129 727
rect -369 655 -353 689
rect -319 655 -303 689
rect -369 639 -303 655
rect -177 689 -111 705
rect -63 701 -33 727
rect 33 705 63 727
rect -177 655 -161 689
rect -127 655 -111 689
rect -177 639 -111 655
rect 15 689 81 705
rect 129 701 159 727
rect 225 705 255 727
rect 15 655 31 689
rect 65 655 81 689
rect 15 639 81 655
rect 207 689 273 705
rect 321 701 351 727
rect 417 705 447 727
rect 207 655 223 689
rect 257 655 273 689
rect 207 639 273 655
rect 399 689 465 705
rect 513 701 543 727
rect 609 705 639 727
rect 399 655 415 689
rect 449 655 465 689
rect 399 639 465 655
rect 591 689 657 705
rect 705 701 735 727
rect 801 705 831 727
rect 591 655 607 689
rect 641 655 657 689
rect 591 639 657 655
rect 783 689 849 705
rect 897 701 927 727
rect 993 705 1023 727
rect 783 655 799 689
rect 833 655 849 689
rect 783 639 849 655
rect 975 689 1041 705
rect 1089 701 1119 727
rect 1185 705 1215 727
rect 975 655 991 689
rect 1025 655 1041 689
rect 975 639 1041 655
rect 1167 689 1233 705
rect 1281 701 1311 727
rect 1377 705 1407 727
rect 1167 655 1183 689
rect 1217 655 1233 689
rect 1167 639 1233 655
rect 1359 689 1425 705
rect 1473 701 1503 727
rect 1569 705 1599 727
rect 1359 655 1375 689
rect 1409 655 1425 689
rect 1359 639 1425 655
rect 1551 689 1617 705
rect 1665 701 1695 727
rect 1761 705 1791 727
rect 1551 655 1567 689
rect 1601 655 1617 689
rect 1551 639 1617 655
rect 1743 689 1809 705
rect 1857 701 1887 727
rect 1953 705 1983 727
rect 1743 655 1759 689
rect 1793 655 1809 689
rect 1743 639 1809 655
rect 1935 689 2001 705
rect 2049 701 2079 727
rect 2145 705 2175 727
rect 1935 655 1951 689
rect 1985 655 2001 689
rect 1935 639 2001 655
rect 2127 689 2193 705
rect 2241 701 2271 727
rect 2337 705 2367 727
rect 2127 655 2143 689
rect 2177 655 2193 689
rect 2127 639 2193 655
rect 2319 689 2385 705
rect 2319 655 2335 689
rect 2369 655 2385 689
rect 2319 639 2385 655
rect -2289 581 -2223 597
rect -2289 547 -2273 581
rect -2239 547 -2223 581
rect -2367 509 -2337 535
rect -2289 531 -2223 547
rect -2097 581 -2031 597
rect -2097 547 -2081 581
rect -2047 547 -2031 581
rect -2271 509 -2241 531
rect -2175 509 -2145 535
rect -2097 531 -2031 547
rect -1905 581 -1839 597
rect -1905 547 -1889 581
rect -1855 547 -1839 581
rect -2079 509 -2049 531
rect -1983 509 -1953 535
rect -1905 531 -1839 547
rect -1713 581 -1647 597
rect -1713 547 -1697 581
rect -1663 547 -1647 581
rect -1887 509 -1857 531
rect -1791 509 -1761 535
rect -1713 531 -1647 547
rect -1521 581 -1455 597
rect -1521 547 -1505 581
rect -1471 547 -1455 581
rect -1695 509 -1665 531
rect -1599 509 -1569 535
rect -1521 531 -1455 547
rect -1329 581 -1263 597
rect -1329 547 -1313 581
rect -1279 547 -1263 581
rect -1503 509 -1473 531
rect -1407 509 -1377 535
rect -1329 531 -1263 547
rect -1137 581 -1071 597
rect -1137 547 -1121 581
rect -1087 547 -1071 581
rect -1311 509 -1281 531
rect -1215 509 -1185 535
rect -1137 531 -1071 547
rect -945 581 -879 597
rect -945 547 -929 581
rect -895 547 -879 581
rect -1119 509 -1089 531
rect -1023 509 -993 535
rect -945 531 -879 547
rect -753 581 -687 597
rect -753 547 -737 581
rect -703 547 -687 581
rect -927 509 -897 531
rect -831 509 -801 535
rect -753 531 -687 547
rect -561 581 -495 597
rect -561 547 -545 581
rect -511 547 -495 581
rect -735 509 -705 531
rect -639 509 -609 535
rect -561 531 -495 547
rect -369 581 -303 597
rect -369 547 -353 581
rect -319 547 -303 581
rect -543 509 -513 531
rect -447 509 -417 535
rect -369 531 -303 547
rect -177 581 -111 597
rect -177 547 -161 581
rect -127 547 -111 581
rect -351 509 -321 531
rect -255 509 -225 535
rect -177 531 -111 547
rect 15 581 81 597
rect 15 547 31 581
rect 65 547 81 581
rect -159 509 -129 531
rect -63 509 -33 535
rect 15 531 81 547
rect 207 581 273 597
rect 207 547 223 581
rect 257 547 273 581
rect 33 509 63 531
rect 129 509 159 535
rect 207 531 273 547
rect 399 581 465 597
rect 399 547 415 581
rect 449 547 465 581
rect 225 509 255 531
rect 321 509 351 535
rect 399 531 465 547
rect 591 581 657 597
rect 591 547 607 581
rect 641 547 657 581
rect 417 509 447 531
rect 513 509 543 535
rect 591 531 657 547
rect 783 581 849 597
rect 783 547 799 581
rect 833 547 849 581
rect 609 509 639 531
rect 705 509 735 535
rect 783 531 849 547
rect 975 581 1041 597
rect 975 547 991 581
rect 1025 547 1041 581
rect 801 509 831 531
rect 897 509 927 535
rect 975 531 1041 547
rect 1167 581 1233 597
rect 1167 547 1183 581
rect 1217 547 1233 581
rect 993 509 1023 531
rect 1089 509 1119 535
rect 1167 531 1233 547
rect 1359 581 1425 597
rect 1359 547 1375 581
rect 1409 547 1425 581
rect 1185 509 1215 531
rect 1281 509 1311 535
rect 1359 531 1425 547
rect 1551 581 1617 597
rect 1551 547 1567 581
rect 1601 547 1617 581
rect 1377 509 1407 531
rect 1473 509 1503 535
rect 1551 531 1617 547
rect 1743 581 1809 597
rect 1743 547 1759 581
rect 1793 547 1809 581
rect 1569 509 1599 531
rect 1665 509 1695 535
rect 1743 531 1809 547
rect 1935 581 2001 597
rect 1935 547 1951 581
rect 1985 547 2001 581
rect 1761 509 1791 531
rect 1857 509 1887 535
rect 1935 531 2001 547
rect 2127 581 2193 597
rect 2127 547 2143 581
rect 2177 547 2193 581
rect 1953 509 1983 531
rect 2049 509 2079 535
rect 2127 531 2193 547
rect 2319 581 2385 597
rect 2319 547 2335 581
rect 2369 547 2385 581
rect 2145 509 2175 531
rect 2241 509 2271 535
rect 2319 531 2385 547
rect 2337 509 2367 531
rect -2367 87 -2337 109
rect -2385 71 -2319 87
rect -2271 83 -2241 109
rect -2175 87 -2145 109
rect -2385 37 -2369 71
rect -2335 37 -2319 71
rect -2385 21 -2319 37
rect -2193 71 -2127 87
rect -2079 83 -2049 109
rect -1983 87 -1953 109
rect -2193 37 -2177 71
rect -2143 37 -2127 71
rect -2193 21 -2127 37
rect -2001 71 -1935 87
rect -1887 83 -1857 109
rect -1791 87 -1761 109
rect -2001 37 -1985 71
rect -1951 37 -1935 71
rect -2001 21 -1935 37
rect -1809 71 -1743 87
rect -1695 83 -1665 109
rect -1599 87 -1569 109
rect -1809 37 -1793 71
rect -1759 37 -1743 71
rect -1809 21 -1743 37
rect -1617 71 -1551 87
rect -1503 83 -1473 109
rect -1407 87 -1377 109
rect -1617 37 -1601 71
rect -1567 37 -1551 71
rect -1617 21 -1551 37
rect -1425 71 -1359 87
rect -1311 83 -1281 109
rect -1215 87 -1185 109
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1425 21 -1359 37
rect -1233 71 -1167 87
rect -1119 83 -1089 109
rect -1023 87 -993 109
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1233 21 -1167 37
rect -1041 71 -975 87
rect -927 83 -897 109
rect -831 87 -801 109
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -1041 21 -975 37
rect -849 71 -783 87
rect -735 83 -705 109
rect -639 87 -609 109
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -543 83 -513 109
rect -447 87 -417 109
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 513 87 543 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 609 83 639 109
rect 705 87 735 109
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 801 83 831 109
rect 897 87 927 109
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 993 83 1023 109
rect 1089 87 1119 109
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect 1071 71 1137 87
rect 1185 83 1215 109
rect 1281 87 1311 109
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1071 21 1137 37
rect 1263 71 1329 87
rect 1377 83 1407 109
rect 1473 87 1503 109
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1263 21 1329 37
rect 1455 71 1521 87
rect 1569 83 1599 109
rect 1665 87 1695 109
rect 1455 37 1471 71
rect 1505 37 1521 71
rect 1455 21 1521 37
rect 1647 71 1713 87
rect 1761 83 1791 109
rect 1857 87 1887 109
rect 1647 37 1663 71
rect 1697 37 1713 71
rect 1647 21 1713 37
rect 1839 71 1905 87
rect 1953 83 1983 109
rect 2049 87 2079 109
rect 1839 37 1855 71
rect 1889 37 1905 71
rect 1839 21 1905 37
rect 2031 71 2097 87
rect 2145 83 2175 109
rect 2241 87 2271 109
rect 2031 37 2047 71
rect 2081 37 2097 71
rect 2031 21 2097 37
rect 2223 71 2289 87
rect 2337 83 2367 109
rect 2223 37 2239 71
rect 2273 37 2289 71
rect 2223 21 2289 37
rect -2385 -37 -2319 -21
rect -2385 -71 -2369 -37
rect -2335 -71 -2319 -37
rect -2385 -87 -2319 -71
rect -2193 -37 -2127 -21
rect -2193 -71 -2177 -37
rect -2143 -71 -2127 -37
rect -2367 -109 -2337 -87
rect -2271 -109 -2241 -83
rect -2193 -87 -2127 -71
rect -2001 -37 -1935 -21
rect -2001 -71 -1985 -37
rect -1951 -71 -1935 -37
rect -2175 -109 -2145 -87
rect -2079 -109 -2049 -83
rect -2001 -87 -1935 -71
rect -1809 -37 -1743 -21
rect -1809 -71 -1793 -37
rect -1759 -71 -1743 -37
rect -1983 -109 -1953 -87
rect -1887 -109 -1857 -83
rect -1809 -87 -1743 -71
rect -1617 -37 -1551 -21
rect -1617 -71 -1601 -37
rect -1567 -71 -1551 -37
rect -1791 -109 -1761 -87
rect -1695 -109 -1665 -83
rect -1617 -87 -1551 -71
rect -1425 -37 -1359 -21
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1599 -109 -1569 -87
rect -1503 -109 -1473 -83
rect -1425 -87 -1359 -71
rect -1233 -37 -1167 -21
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1407 -109 -1377 -87
rect -1311 -109 -1281 -83
rect -1233 -87 -1167 -71
rect -1041 -37 -975 -21
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -1215 -109 -1185 -87
rect -1119 -109 -1089 -83
rect -1041 -87 -975 -71
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -1023 -109 -993 -87
rect -927 -109 -897 -83
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -831 -109 -801 -87
rect -735 -109 -705 -83
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -639 -109 -609 -87
rect -543 -109 -513 -83
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 321 -109 351 -87
rect 417 -109 447 -83
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 513 -109 543 -87
rect 609 -109 639 -83
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 705 -109 735 -87
rect 801 -109 831 -83
rect 879 -87 945 -71
rect 1071 -37 1137 -21
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 897 -109 927 -87
rect 993 -109 1023 -83
rect 1071 -87 1137 -71
rect 1263 -37 1329 -21
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1089 -109 1119 -87
rect 1185 -109 1215 -83
rect 1263 -87 1329 -71
rect 1455 -37 1521 -21
rect 1455 -71 1471 -37
rect 1505 -71 1521 -37
rect 1281 -109 1311 -87
rect 1377 -109 1407 -83
rect 1455 -87 1521 -71
rect 1647 -37 1713 -21
rect 1647 -71 1663 -37
rect 1697 -71 1713 -37
rect 1473 -109 1503 -87
rect 1569 -109 1599 -83
rect 1647 -87 1713 -71
rect 1839 -37 1905 -21
rect 1839 -71 1855 -37
rect 1889 -71 1905 -37
rect 1665 -109 1695 -87
rect 1761 -109 1791 -83
rect 1839 -87 1905 -71
rect 2031 -37 2097 -21
rect 2031 -71 2047 -37
rect 2081 -71 2097 -37
rect 1857 -109 1887 -87
rect 1953 -109 1983 -83
rect 2031 -87 2097 -71
rect 2223 -37 2289 -21
rect 2223 -71 2239 -37
rect 2273 -71 2289 -37
rect 2049 -109 2079 -87
rect 2145 -109 2175 -83
rect 2223 -87 2289 -71
rect 2241 -109 2271 -87
rect 2337 -109 2367 -83
rect -2367 -535 -2337 -509
rect -2271 -531 -2241 -509
rect -2289 -547 -2223 -531
rect -2175 -535 -2145 -509
rect -2079 -531 -2049 -509
rect -2289 -581 -2273 -547
rect -2239 -581 -2223 -547
rect -2289 -597 -2223 -581
rect -2097 -547 -2031 -531
rect -1983 -535 -1953 -509
rect -1887 -531 -1857 -509
rect -2097 -581 -2081 -547
rect -2047 -581 -2031 -547
rect -2097 -597 -2031 -581
rect -1905 -547 -1839 -531
rect -1791 -535 -1761 -509
rect -1695 -531 -1665 -509
rect -1905 -581 -1889 -547
rect -1855 -581 -1839 -547
rect -1905 -597 -1839 -581
rect -1713 -547 -1647 -531
rect -1599 -535 -1569 -509
rect -1503 -531 -1473 -509
rect -1713 -581 -1697 -547
rect -1663 -581 -1647 -547
rect -1713 -597 -1647 -581
rect -1521 -547 -1455 -531
rect -1407 -535 -1377 -509
rect -1311 -531 -1281 -509
rect -1521 -581 -1505 -547
rect -1471 -581 -1455 -547
rect -1521 -597 -1455 -581
rect -1329 -547 -1263 -531
rect -1215 -535 -1185 -509
rect -1119 -531 -1089 -509
rect -1329 -581 -1313 -547
rect -1279 -581 -1263 -547
rect -1329 -597 -1263 -581
rect -1137 -547 -1071 -531
rect -1023 -535 -993 -509
rect -927 -531 -897 -509
rect -1137 -581 -1121 -547
rect -1087 -581 -1071 -547
rect -1137 -597 -1071 -581
rect -945 -547 -879 -531
rect -831 -535 -801 -509
rect -735 -531 -705 -509
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -945 -597 -879 -581
rect -753 -547 -687 -531
rect -639 -535 -609 -509
rect -543 -531 -513 -509
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -753 -597 -687 -581
rect -561 -547 -495 -531
rect -447 -535 -417 -509
rect -351 -531 -321 -509
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -561 -597 -495 -581
rect -369 -547 -303 -531
rect -255 -535 -225 -509
rect -159 -531 -129 -509
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -369 -597 -303 -581
rect -177 -547 -111 -531
rect -63 -535 -33 -509
rect 33 -531 63 -509
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 129 -535 159 -509
rect 225 -531 255 -509
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
rect 207 -547 273 -531
rect 321 -535 351 -509
rect 417 -531 447 -509
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 207 -597 273 -581
rect 399 -547 465 -531
rect 513 -535 543 -509
rect 609 -531 639 -509
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 399 -597 465 -581
rect 591 -547 657 -531
rect 705 -535 735 -509
rect 801 -531 831 -509
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 591 -597 657 -581
rect 783 -547 849 -531
rect 897 -535 927 -509
rect 993 -531 1023 -509
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 783 -597 849 -581
rect 975 -547 1041 -531
rect 1089 -535 1119 -509
rect 1185 -531 1215 -509
rect 975 -581 991 -547
rect 1025 -581 1041 -547
rect 975 -597 1041 -581
rect 1167 -547 1233 -531
rect 1281 -535 1311 -509
rect 1377 -531 1407 -509
rect 1167 -581 1183 -547
rect 1217 -581 1233 -547
rect 1167 -597 1233 -581
rect 1359 -547 1425 -531
rect 1473 -535 1503 -509
rect 1569 -531 1599 -509
rect 1359 -581 1375 -547
rect 1409 -581 1425 -547
rect 1359 -597 1425 -581
rect 1551 -547 1617 -531
rect 1665 -535 1695 -509
rect 1761 -531 1791 -509
rect 1551 -581 1567 -547
rect 1601 -581 1617 -547
rect 1551 -597 1617 -581
rect 1743 -547 1809 -531
rect 1857 -535 1887 -509
rect 1953 -531 1983 -509
rect 1743 -581 1759 -547
rect 1793 -581 1809 -547
rect 1743 -597 1809 -581
rect 1935 -547 2001 -531
rect 2049 -535 2079 -509
rect 2145 -531 2175 -509
rect 1935 -581 1951 -547
rect 1985 -581 2001 -547
rect 1935 -597 2001 -581
rect 2127 -547 2193 -531
rect 2241 -535 2271 -509
rect 2337 -531 2367 -509
rect 2127 -581 2143 -547
rect 2177 -581 2193 -547
rect 2127 -597 2193 -581
rect 2319 -547 2385 -531
rect 2319 -581 2335 -547
rect 2369 -581 2385 -547
rect 2319 -597 2385 -581
rect -2289 -655 -2223 -639
rect -2289 -689 -2273 -655
rect -2239 -689 -2223 -655
rect -2367 -727 -2337 -701
rect -2289 -705 -2223 -689
rect -2097 -655 -2031 -639
rect -2097 -689 -2081 -655
rect -2047 -689 -2031 -655
rect -2271 -727 -2241 -705
rect -2175 -727 -2145 -701
rect -2097 -705 -2031 -689
rect -1905 -655 -1839 -639
rect -1905 -689 -1889 -655
rect -1855 -689 -1839 -655
rect -2079 -727 -2049 -705
rect -1983 -727 -1953 -701
rect -1905 -705 -1839 -689
rect -1713 -655 -1647 -639
rect -1713 -689 -1697 -655
rect -1663 -689 -1647 -655
rect -1887 -727 -1857 -705
rect -1791 -727 -1761 -701
rect -1713 -705 -1647 -689
rect -1521 -655 -1455 -639
rect -1521 -689 -1505 -655
rect -1471 -689 -1455 -655
rect -1695 -727 -1665 -705
rect -1599 -727 -1569 -701
rect -1521 -705 -1455 -689
rect -1329 -655 -1263 -639
rect -1329 -689 -1313 -655
rect -1279 -689 -1263 -655
rect -1503 -727 -1473 -705
rect -1407 -727 -1377 -701
rect -1329 -705 -1263 -689
rect -1137 -655 -1071 -639
rect -1137 -689 -1121 -655
rect -1087 -689 -1071 -655
rect -1311 -727 -1281 -705
rect -1215 -727 -1185 -701
rect -1137 -705 -1071 -689
rect -945 -655 -879 -639
rect -945 -689 -929 -655
rect -895 -689 -879 -655
rect -1119 -727 -1089 -705
rect -1023 -727 -993 -701
rect -945 -705 -879 -689
rect -753 -655 -687 -639
rect -753 -689 -737 -655
rect -703 -689 -687 -655
rect -927 -727 -897 -705
rect -831 -727 -801 -701
rect -753 -705 -687 -689
rect -561 -655 -495 -639
rect -561 -689 -545 -655
rect -511 -689 -495 -655
rect -735 -727 -705 -705
rect -639 -727 -609 -701
rect -561 -705 -495 -689
rect -369 -655 -303 -639
rect -369 -689 -353 -655
rect -319 -689 -303 -655
rect -543 -727 -513 -705
rect -447 -727 -417 -701
rect -369 -705 -303 -689
rect -177 -655 -111 -639
rect -177 -689 -161 -655
rect -127 -689 -111 -655
rect -351 -727 -321 -705
rect -255 -727 -225 -701
rect -177 -705 -111 -689
rect 15 -655 81 -639
rect 15 -689 31 -655
rect 65 -689 81 -655
rect -159 -727 -129 -705
rect -63 -727 -33 -701
rect 15 -705 81 -689
rect 207 -655 273 -639
rect 207 -689 223 -655
rect 257 -689 273 -655
rect 33 -727 63 -705
rect 129 -727 159 -701
rect 207 -705 273 -689
rect 399 -655 465 -639
rect 399 -689 415 -655
rect 449 -689 465 -655
rect 225 -727 255 -705
rect 321 -727 351 -701
rect 399 -705 465 -689
rect 591 -655 657 -639
rect 591 -689 607 -655
rect 641 -689 657 -655
rect 417 -727 447 -705
rect 513 -727 543 -701
rect 591 -705 657 -689
rect 783 -655 849 -639
rect 783 -689 799 -655
rect 833 -689 849 -655
rect 609 -727 639 -705
rect 705 -727 735 -701
rect 783 -705 849 -689
rect 975 -655 1041 -639
rect 975 -689 991 -655
rect 1025 -689 1041 -655
rect 801 -727 831 -705
rect 897 -727 927 -701
rect 975 -705 1041 -689
rect 1167 -655 1233 -639
rect 1167 -689 1183 -655
rect 1217 -689 1233 -655
rect 993 -727 1023 -705
rect 1089 -727 1119 -701
rect 1167 -705 1233 -689
rect 1359 -655 1425 -639
rect 1359 -689 1375 -655
rect 1409 -689 1425 -655
rect 1185 -727 1215 -705
rect 1281 -727 1311 -701
rect 1359 -705 1425 -689
rect 1551 -655 1617 -639
rect 1551 -689 1567 -655
rect 1601 -689 1617 -655
rect 1377 -727 1407 -705
rect 1473 -727 1503 -701
rect 1551 -705 1617 -689
rect 1743 -655 1809 -639
rect 1743 -689 1759 -655
rect 1793 -689 1809 -655
rect 1569 -727 1599 -705
rect 1665 -727 1695 -701
rect 1743 -705 1809 -689
rect 1935 -655 2001 -639
rect 1935 -689 1951 -655
rect 1985 -689 2001 -655
rect 1761 -727 1791 -705
rect 1857 -727 1887 -701
rect 1935 -705 2001 -689
rect 2127 -655 2193 -639
rect 2127 -689 2143 -655
rect 2177 -689 2193 -655
rect 1953 -727 1983 -705
rect 2049 -727 2079 -701
rect 2127 -705 2193 -689
rect 2319 -655 2385 -639
rect 2319 -689 2335 -655
rect 2369 -689 2385 -655
rect 2145 -727 2175 -705
rect 2241 -727 2271 -701
rect 2319 -705 2385 -689
rect 2337 -727 2367 -705
rect -2367 -1149 -2337 -1127
rect -2385 -1165 -2319 -1149
rect -2271 -1153 -2241 -1127
rect -2175 -1149 -2145 -1127
rect -2385 -1199 -2369 -1165
rect -2335 -1199 -2319 -1165
rect -2385 -1215 -2319 -1199
rect -2193 -1165 -2127 -1149
rect -2079 -1153 -2049 -1127
rect -1983 -1149 -1953 -1127
rect -2193 -1199 -2177 -1165
rect -2143 -1199 -2127 -1165
rect -2193 -1215 -2127 -1199
rect -2001 -1165 -1935 -1149
rect -1887 -1153 -1857 -1127
rect -1791 -1149 -1761 -1127
rect -2001 -1199 -1985 -1165
rect -1951 -1199 -1935 -1165
rect -2001 -1215 -1935 -1199
rect -1809 -1165 -1743 -1149
rect -1695 -1153 -1665 -1127
rect -1599 -1149 -1569 -1127
rect -1809 -1199 -1793 -1165
rect -1759 -1199 -1743 -1165
rect -1809 -1215 -1743 -1199
rect -1617 -1165 -1551 -1149
rect -1503 -1153 -1473 -1127
rect -1407 -1149 -1377 -1127
rect -1617 -1199 -1601 -1165
rect -1567 -1199 -1551 -1165
rect -1617 -1215 -1551 -1199
rect -1425 -1165 -1359 -1149
rect -1311 -1153 -1281 -1127
rect -1215 -1149 -1185 -1127
rect -1425 -1199 -1409 -1165
rect -1375 -1199 -1359 -1165
rect -1425 -1215 -1359 -1199
rect -1233 -1165 -1167 -1149
rect -1119 -1153 -1089 -1127
rect -1023 -1149 -993 -1127
rect -1233 -1199 -1217 -1165
rect -1183 -1199 -1167 -1165
rect -1233 -1215 -1167 -1199
rect -1041 -1165 -975 -1149
rect -927 -1153 -897 -1127
rect -831 -1149 -801 -1127
rect -1041 -1199 -1025 -1165
rect -991 -1199 -975 -1165
rect -1041 -1215 -975 -1199
rect -849 -1165 -783 -1149
rect -735 -1153 -705 -1127
rect -639 -1149 -609 -1127
rect -849 -1199 -833 -1165
rect -799 -1199 -783 -1165
rect -849 -1215 -783 -1199
rect -657 -1165 -591 -1149
rect -543 -1153 -513 -1127
rect -447 -1149 -417 -1127
rect -657 -1199 -641 -1165
rect -607 -1199 -591 -1165
rect -657 -1215 -591 -1199
rect -465 -1165 -399 -1149
rect -351 -1153 -321 -1127
rect -255 -1149 -225 -1127
rect -465 -1199 -449 -1165
rect -415 -1199 -399 -1165
rect -465 -1215 -399 -1199
rect -273 -1165 -207 -1149
rect -159 -1153 -129 -1127
rect -63 -1149 -33 -1127
rect -273 -1199 -257 -1165
rect -223 -1199 -207 -1165
rect -273 -1215 -207 -1199
rect -81 -1165 -15 -1149
rect 33 -1153 63 -1127
rect 129 -1149 159 -1127
rect -81 -1199 -65 -1165
rect -31 -1199 -15 -1165
rect -81 -1215 -15 -1199
rect 111 -1165 177 -1149
rect 225 -1153 255 -1127
rect 321 -1149 351 -1127
rect 111 -1199 127 -1165
rect 161 -1199 177 -1165
rect 111 -1215 177 -1199
rect 303 -1165 369 -1149
rect 417 -1153 447 -1127
rect 513 -1149 543 -1127
rect 303 -1199 319 -1165
rect 353 -1199 369 -1165
rect 303 -1215 369 -1199
rect 495 -1165 561 -1149
rect 609 -1153 639 -1127
rect 705 -1149 735 -1127
rect 495 -1199 511 -1165
rect 545 -1199 561 -1165
rect 495 -1215 561 -1199
rect 687 -1165 753 -1149
rect 801 -1153 831 -1127
rect 897 -1149 927 -1127
rect 687 -1199 703 -1165
rect 737 -1199 753 -1165
rect 687 -1215 753 -1199
rect 879 -1165 945 -1149
rect 993 -1153 1023 -1127
rect 1089 -1149 1119 -1127
rect 879 -1199 895 -1165
rect 929 -1199 945 -1165
rect 879 -1215 945 -1199
rect 1071 -1165 1137 -1149
rect 1185 -1153 1215 -1127
rect 1281 -1149 1311 -1127
rect 1071 -1199 1087 -1165
rect 1121 -1199 1137 -1165
rect 1071 -1215 1137 -1199
rect 1263 -1165 1329 -1149
rect 1377 -1153 1407 -1127
rect 1473 -1149 1503 -1127
rect 1263 -1199 1279 -1165
rect 1313 -1199 1329 -1165
rect 1263 -1215 1329 -1199
rect 1455 -1165 1521 -1149
rect 1569 -1153 1599 -1127
rect 1665 -1149 1695 -1127
rect 1455 -1199 1471 -1165
rect 1505 -1199 1521 -1165
rect 1455 -1215 1521 -1199
rect 1647 -1165 1713 -1149
rect 1761 -1153 1791 -1127
rect 1857 -1149 1887 -1127
rect 1647 -1199 1663 -1165
rect 1697 -1199 1713 -1165
rect 1647 -1215 1713 -1199
rect 1839 -1165 1905 -1149
rect 1953 -1153 1983 -1127
rect 2049 -1149 2079 -1127
rect 1839 -1199 1855 -1165
rect 1889 -1199 1905 -1165
rect 1839 -1215 1905 -1199
rect 2031 -1165 2097 -1149
rect 2145 -1153 2175 -1127
rect 2241 -1149 2271 -1127
rect 2031 -1199 2047 -1165
rect 2081 -1199 2097 -1165
rect 2031 -1215 2097 -1199
rect 2223 -1165 2289 -1149
rect 2337 -1153 2367 -1127
rect 2223 -1199 2239 -1165
rect 2273 -1199 2289 -1165
rect 2223 -1215 2289 -1199
<< polycont >>
rect -2369 1165 -2335 1199
rect -2177 1165 -2143 1199
rect -1985 1165 -1951 1199
rect -1793 1165 -1759 1199
rect -1601 1165 -1567 1199
rect -1409 1165 -1375 1199
rect -1217 1165 -1183 1199
rect -1025 1165 -991 1199
rect -833 1165 -799 1199
rect -641 1165 -607 1199
rect -449 1165 -415 1199
rect -257 1165 -223 1199
rect -65 1165 -31 1199
rect 127 1165 161 1199
rect 319 1165 353 1199
rect 511 1165 545 1199
rect 703 1165 737 1199
rect 895 1165 929 1199
rect 1087 1165 1121 1199
rect 1279 1165 1313 1199
rect 1471 1165 1505 1199
rect 1663 1165 1697 1199
rect 1855 1165 1889 1199
rect 2047 1165 2081 1199
rect 2239 1165 2273 1199
rect -2273 655 -2239 689
rect -2081 655 -2047 689
rect -1889 655 -1855 689
rect -1697 655 -1663 689
rect -1505 655 -1471 689
rect -1313 655 -1279 689
rect -1121 655 -1087 689
rect -929 655 -895 689
rect -737 655 -703 689
rect -545 655 -511 689
rect -353 655 -319 689
rect -161 655 -127 689
rect 31 655 65 689
rect 223 655 257 689
rect 415 655 449 689
rect 607 655 641 689
rect 799 655 833 689
rect 991 655 1025 689
rect 1183 655 1217 689
rect 1375 655 1409 689
rect 1567 655 1601 689
rect 1759 655 1793 689
rect 1951 655 1985 689
rect 2143 655 2177 689
rect 2335 655 2369 689
rect -2273 547 -2239 581
rect -2081 547 -2047 581
rect -1889 547 -1855 581
rect -1697 547 -1663 581
rect -1505 547 -1471 581
rect -1313 547 -1279 581
rect -1121 547 -1087 581
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect 991 547 1025 581
rect 1183 547 1217 581
rect 1375 547 1409 581
rect 1567 547 1601 581
rect 1759 547 1793 581
rect 1951 547 1985 581
rect 2143 547 2177 581
rect 2335 547 2369 581
rect -2369 37 -2335 71
rect -2177 37 -2143 71
rect -1985 37 -1951 71
rect -1793 37 -1759 71
rect -1601 37 -1567 71
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect 1471 37 1505 71
rect 1663 37 1697 71
rect 1855 37 1889 71
rect 2047 37 2081 71
rect 2239 37 2273 71
rect -2369 -71 -2335 -37
rect -2177 -71 -2143 -37
rect -1985 -71 -1951 -37
rect -1793 -71 -1759 -37
rect -1601 -71 -1567 -37
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect 1471 -71 1505 -37
rect 1663 -71 1697 -37
rect 1855 -71 1889 -37
rect 2047 -71 2081 -37
rect 2239 -71 2273 -37
rect -2273 -581 -2239 -547
rect -2081 -581 -2047 -547
rect -1889 -581 -1855 -547
rect -1697 -581 -1663 -547
rect -1505 -581 -1471 -547
rect -1313 -581 -1279 -547
rect -1121 -581 -1087 -547
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
rect 991 -581 1025 -547
rect 1183 -581 1217 -547
rect 1375 -581 1409 -547
rect 1567 -581 1601 -547
rect 1759 -581 1793 -547
rect 1951 -581 1985 -547
rect 2143 -581 2177 -547
rect 2335 -581 2369 -547
rect -2273 -689 -2239 -655
rect -2081 -689 -2047 -655
rect -1889 -689 -1855 -655
rect -1697 -689 -1663 -655
rect -1505 -689 -1471 -655
rect -1313 -689 -1279 -655
rect -1121 -689 -1087 -655
rect -929 -689 -895 -655
rect -737 -689 -703 -655
rect -545 -689 -511 -655
rect -353 -689 -319 -655
rect -161 -689 -127 -655
rect 31 -689 65 -655
rect 223 -689 257 -655
rect 415 -689 449 -655
rect 607 -689 641 -655
rect 799 -689 833 -655
rect 991 -689 1025 -655
rect 1183 -689 1217 -655
rect 1375 -689 1409 -655
rect 1567 -689 1601 -655
rect 1759 -689 1793 -655
rect 1951 -689 1985 -655
rect 2143 -689 2177 -655
rect 2335 -689 2369 -655
rect -2369 -1199 -2335 -1165
rect -2177 -1199 -2143 -1165
rect -1985 -1199 -1951 -1165
rect -1793 -1199 -1759 -1165
rect -1601 -1199 -1567 -1165
rect -1409 -1199 -1375 -1165
rect -1217 -1199 -1183 -1165
rect -1025 -1199 -991 -1165
rect -833 -1199 -799 -1165
rect -641 -1199 -607 -1165
rect -449 -1199 -415 -1165
rect -257 -1199 -223 -1165
rect -65 -1199 -31 -1165
rect 127 -1199 161 -1165
rect 319 -1199 353 -1165
rect 511 -1199 545 -1165
rect 703 -1199 737 -1165
rect 895 -1199 929 -1165
rect 1087 -1199 1121 -1165
rect 1279 -1199 1313 -1165
rect 1471 -1199 1505 -1165
rect 1663 -1199 1697 -1165
rect 1855 -1199 1889 -1165
rect 2047 -1199 2081 -1165
rect 2239 -1199 2273 -1165
<< locali >>
rect -2531 1267 -2435 1301
rect 2435 1267 2531 1301
rect -2531 1205 -2497 1267
rect 2497 1205 2531 1267
rect -2385 1165 -2369 1199
rect -2335 1165 -2319 1199
rect -2193 1165 -2177 1199
rect -2143 1165 -2127 1199
rect -2001 1165 -1985 1199
rect -1951 1165 -1935 1199
rect -1809 1165 -1793 1199
rect -1759 1165 -1743 1199
rect -1617 1165 -1601 1199
rect -1567 1165 -1551 1199
rect -1425 1165 -1409 1199
rect -1375 1165 -1359 1199
rect -1233 1165 -1217 1199
rect -1183 1165 -1167 1199
rect -1041 1165 -1025 1199
rect -991 1165 -975 1199
rect -849 1165 -833 1199
rect -799 1165 -783 1199
rect -657 1165 -641 1199
rect -607 1165 -591 1199
rect -465 1165 -449 1199
rect -415 1165 -399 1199
rect -273 1165 -257 1199
rect -223 1165 -207 1199
rect -81 1165 -65 1199
rect -31 1165 -15 1199
rect 111 1165 127 1199
rect 161 1165 177 1199
rect 303 1165 319 1199
rect 353 1165 369 1199
rect 495 1165 511 1199
rect 545 1165 561 1199
rect 687 1165 703 1199
rect 737 1165 753 1199
rect 879 1165 895 1199
rect 929 1165 945 1199
rect 1071 1165 1087 1199
rect 1121 1165 1137 1199
rect 1263 1165 1279 1199
rect 1313 1165 1329 1199
rect 1455 1165 1471 1199
rect 1505 1165 1521 1199
rect 1647 1165 1663 1199
rect 1697 1165 1713 1199
rect 1839 1165 1855 1199
rect 1889 1165 1905 1199
rect 2031 1165 2047 1199
rect 2081 1165 2097 1199
rect 2223 1165 2239 1199
rect 2273 1165 2289 1199
rect -2417 1115 -2383 1131
rect -2417 723 -2383 739
rect -2321 1115 -2287 1131
rect -2321 723 -2287 739
rect -2225 1115 -2191 1131
rect -2225 723 -2191 739
rect -2129 1115 -2095 1131
rect -2129 723 -2095 739
rect -2033 1115 -1999 1131
rect -2033 723 -1999 739
rect -1937 1115 -1903 1131
rect -1937 723 -1903 739
rect -1841 1115 -1807 1131
rect -1841 723 -1807 739
rect -1745 1115 -1711 1131
rect -1745 723 -1711 739
rect -1649 1115 -1615 1131
rect -1649 723 -1615 739
rect -1553 1115 -1519 1131
rect -1553 723 -1519 739
rect -1457 1115 -1423 1131
rect -1457 723 -1423 739
rect -1361 1115 -1327 1131
rect -1361 723 -1327 739
rect -1265 1115 -1231 1131
rect -1265 723 -1231 739
rect -1169 1115 -1135 1131
rect -1169 723 -1135 739
rect -1073 1115 -1039 1131
rect -1073 723 -1039 739
rect -977 1115 -943 1131
rect -977 723 -943 739
rect -881 1115 -847 1131
rect -881 723 -847 739
rect -785 1115 -751 1131
rect -785 723 -751 739
rect -689 1115 -655 1131
rect -689 723 -655 739
rect -593 1115 -559 1131
rect -593 723 -559 739
rect -497 1115 -463 1131
rect -497 723 -463 739
rect -401 1115 -367 1131
rect -401 723 -367 739
rect -305 1115 -271 1131
rect -305 723 -271 739
rect -209 1115 -175 1131
rect -209 723 -175 739
rect -113 1115 -79 1131
rect -113 723 -79 739
rect -17 1115 17 1131
rect -17 723 17 739
rect 79 1115 113 1131
rect 79 723 113 739
rect 175 1115 209 1131
rect 175 723 209 739
rect 271 1115 305 1131
rect 271 723 305 739
rect 367 1115 401 1131
rect 367 723 401 739
rect 463 1115 497 1131
rect 463 723 497 739
rect 559 1115 593 1131
rect 559 723 593 739
rect 655 1115 689 1131
rect 655 723 689 739
rect 751 1115 785 1131
rect 751 723 785 739
rect 847 1115 881 1131
rect 847 723 881 739
rect 943 1115 977 1131
rect 943 723 977 739
rect 1039 1115 1073 1131
rect 1039 723 1073 739
rect 1135 1115 1169 1131
rect 1135 723 1169 739
rect 1231 1115 1265 1131
rect 1231 723 1265 739
rect 1327 1115 1361 1131
rect 1327 723 1361 739
rect 1423 1115 1457 1131
rect 1423 723 1457 739
rect 1519 1115 1553 1131
rect 1519 723 1553 739
rect 1615 1115 1649 1131
rect 1615 723 1649 739
rect 1711 1115 1745 1131
rect 1711 723 1745 739
rect 1807 1115 1841 1131
rect 1807 723 1841 739
rect 1903 1115 1937 1131
rect 1903 723 1937 739
rect 1999 1115 2033 1131
rect 1999 723 2033 739
rect 2095 1115 2129 1131
rect 2095 723 2129 739
rect 2191 1115 2225 1131
rect 2191 723 2225 739
rect 2287 1115 2321 1131
rect 2287 723 2321 739
rect 2383 1115 2417 1131
rect 2383 723 2417 739
rect -2289 655 -2273 689
rect -2239 655 -2223 689
rect -2097 655 -2081 689
rect -2047 655 -2031 689
rect -1905 655 -1889 689
rect -1855 655 -1839 689
rect -1713 655 -1697 689
rect -1663 655 -1647 689
rect -1521 655 -1505 689
rect -1471 655 -1455 689
rect -1329 655 -1313 689
rect -1279 655 -1263 689
rect -1137 655 -1121 689
rect -1087 655 -1071 689
rect -945 655 -929 689
rect -895 655 -879 689
rect -753 655 -737 689
rect -703 655 -687 689
rect -561 655 -545 689
rect -511 655 -495 689
rect -369 655 -353 689
rect -319 655 -303 689
rect -177 655 -161 689
rect -127 655 -111 689
rect 15 655 31 689
rect 65 655 81 689
rect 207 655 223 689
rect 257 655 273 689
rect 399 655 415 689
rect 449 655 465 689
rect 591 655 607 689
rect 641 655 657 689
rect 783 655 799 689
rect 833 655 849 689
rect 975 655 991 689
rect 1025 655 1041 689
rect 1167 655 1183 689
rect 1217 655 1233 689
rect 1359 655 1375 689
rect 1409 655 1425 689
rect 1551 655 1567 689
rect 1601 655 1617 689
rect 1743 655 1759 689
rect 1793 655 1809 689
rect 1935 655 1951 689
rect 1985 655 2001 689
rect 2127 655 2143 689
rect 2177 655 2193 689
rect 2319 655 2335 689
rect 2369 655 2385 689
rect -2289 547 -2273 581
rect -2239 547 -2223 581
rect -2097 547 -2081 581
rect -2047 547 -2031 581
rect -1905 547 -1889 581
rect -1855 547 -1839 581
rect -1713 547 -1697 581
rect -1663 547 -1647 581
rect -1521 547 -1505 581
rect -1471 547 -1455 581
rect -1329 547 -1313 581
rect -1279 547 -1263 581
rect -1137 547 -1121 581
rect -1087 547 -1071 581
rect -945 547 -929 581
rect -895 547 -879 581
rect -753 547 -737 581
rect -703 547 -687 581
rect -561 547 -545 581
rect -511 547 -495 581
rect -369 547 -353 581
rect -319 547 -303 581
rect -177 547 -161 581
rect -127 547 -111 581
rect 15 547 31 581
rect 65 547 81 581
rect 207 547 223 581
rect 257 547 273 581
rect 399 547 415 581
rect 449 547 465 581
rect 591 547 607 581
rect 641 547 657 581
rect 783 547 799 581
rect 833 547 849 581
rect 975 547 991 581
rect 1025 547 1041 581
rect 1167 547 1183 581
rect 1217 547 1233 581
rect 1359 547 1375 581
rect 1409 547 1425 581
rect 1551 547 1567 581
rect 1601 547 1617 581
rect 1743 547 1759 581
rect 1793 547 1809 581
rect 1935 547 1951 581
rect 1985 547 2001 581
rect 2127 547 2143 581
rect 2177 547 2193 581
rect 2319 547 2335 581
rect 2369 547 2385 581
rect -2417 497 -2383 513
rect -2417 105 -2383 121
rect -2321 497 -2287 513
rect -2321 105 -2287 121
rect -2225 497 -2191 513
rect -2225 105 -2191 121
rect -2129 497 -2095 513
rect -2129 105 -2095 121
rect -2033 497 -1999 513
rect -2033 105 -1999 121
rect -1937 497 -1903 513
rect -1937 105 -1903 121
rect -1841 497 -1807 513
rect -1841 105 -1807 121
rect -1745 497 -1711 513
rect -1745 105 -1711 121
rect -1649 497 -1615 513
rect -1649 105 -1615 121
rect -1553 497 -1519 513
rect -1553 105 -1519 121
rect -1457 497 -1423 513
rect -1457 105 -1423 121
rect -1361 497 -1327 513
rect -1361 105 -1327 121
rect -1265 497 -1231 513
rect -1265 105 -1231 121
rect -1169 497 -1135 513
rect -1169 105 -1135 121
rect -1073 497 -1039 513
rect -1073 105 -1039 121
rect -977 497 -943 513
rect -977 105 -943 121
rect -881 497 -847 513
rect -881 105 -847 121
rect -785 497 -751 513
rect -785 105 -751 121
rect -689 497 -655 513
rect -689 105 -655 121
rect -593 497 -559 513
rect -593 105 -559 121
rect -497 497 -463 513
rect -497 105 -463 121
rect -401 497 -367 513
rect -401 105 -367 121
rect -305 497 -271 513
rect -305 105 -271 121
rect -209 497 -175 513
rect -209 105 -175 121
rect -113 497 -79 513
rect -113 105 -79 121
rect -17 497 17 513
rect -17 105 17 121
rect 79 497 113 513
rect 79 105 113 121
rect 175 497 209 513
rect 175 105 209 121
rect 271 497 305 513
rect 271 105 305 121
rect 367 497 401 513
rect 367 105 401 121
rect 463 497 497 513
rect 463 105 497 121
rect 559 497 593 513
rect 559 105 593 121
rect 655 497 689 513
rect 655 105 689 121
rect 751 497 785 513
rect 751 105 785 121
rect 847 497 881 513
rect 847 105 881 121
rect 943 497 977 513
rect 943 105 977 121
rect 1039 497 1073 513
rect 1039 105 1073 121
rect 1135 497 1169 513
rect 1135 105 1169 121
rect 1231 497 1265 513
rect 1231 105 1265 121
rect 1327 497 1361 513
rect 1327 105 1361 121
rect 1423 497 1457 513
rect 1423 105 1457 121
rect 1519 497 1553 513
rect 1519 105 1553 121
rect 1615 497 1649 513
rect 1615 105 1649 121
rect 1711 497 1745 513
rect 1711 105 1745 121
rect 1807 497 1841 513
rect 1807 105 1841 121
rect 1903 497 1937 513
rect 1903 105 1937 121
rect 1999 497 2033 513
rect 1999 105 2033 121
rect 2095 497 2129 513
rect 2095 105 2129 121
rect 2191 497 2225 513
rect 2191 105 2225 121
rect 2287 497 2321 513
rect 2287 105 2321 121
rect 2383 497 2417 513
rect 2383 105 2417 121
rect -2385 37 -2369 71
rect -2335 37 -2319 71
rect -2193 37 -2177 71
rect -2143 37 -2127 71
rect -2001 37 -1985 71
rect -1951 37 -1935 71
rect -1809 37 -1793 71
rect -1759 37 -1743 71
rect -1617 37 -1601 71
rect -1567 37 -1551 71
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1455 37 1471 71
rect 1505 37 1521 71
rect 1647 37 1663 71
rect 1697 37 1713 71
rect 1839 37 1855 71
rect 1889 37 1905 71
rect 2031 37 2047 71
rect 2081 37 2097 71
rect 2223 37 2239 71
rect 2273 37 2289 71
rect -2385 -71 -2369 -37
rect -2335 -71 -2319 -37
rect -2193 -71 -2177 -37
rect -2143 -71 -2127 -37
rect -2001 -71 -1985 -37
rect -1951 -71 -1935 -37
rect -1809 -71 -1793 -37
rect -1759 -71 -1743 -37
rect -1617 -71 -1601 -37
rect -1567 -71 -1551 -37
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1455 -71 1471 -37
rect 1505 -71 1521 -37
rect 1647 -71 1663 -37
rect 1697 -71 1713 -37
rect 1839 -71 1855 -37
rect 1889 -71 1905 -37
rect 2031 -71 2047 -37
rect 2081 -71 2097 -37
rect 2223 -71 2239 -37
rect 2273 -71 2289 -37
rect -2417 -121 -2383 -105
rect -2417 -513 -2383 -497
rect -2321 -121 -2287 -105
rect -2321 -513 -2287 -497
rect -2225 -121 -2191 -105
rect -2225 -513 -2191 -497
rect -2129 -121 -2095 -105
rect -2129 -513 -2095 -497
rect -2033 -121 -1999 -105
rect -2033 -513 -1999 -497
rect -1937 -121 -1903 -105
rect -1937 -513 -1903 -497
rect -1841 -121 -1807 -105
rect -1841 -513 -1807 -497
rect -1745 -121 -1711 -105
rect -1745 -513 -1711 -497
rect -1649 -121 -1615 -105
rect -1649 -513 -1615 -497
rect -1553 -121 -1519 -105
rect -1553 -513 -1519 -497
rect -1457 -121 -1423 -105
rect -1457 -513 -1423 -497
rect -1361 -121 -1327 -105
rect -1361 -513 -1327 -497
rect -1265 -121 -1231 -105
rect -1265 -513 -1231 -497
rect -1169 -121 -1135 -105
rect -1169 -513 -1135 -497
rect -1073 -121 -1039 -105
rect -1073 -513 -1039 -497
rect -977 -121 -943 -105
rect -977 -513 -943 -497
rect -881 -121 -847 -105
rect -881 -513 -847 -497
rect -785 -121 -751 -105
rect -785 -513 -751 -497
rect -689 -121 -655 -105
rect -689 -513 -655 -497
rect -593 -121 -559 -105
rect -593 -513 -559 -497
rect -497 -121 -463 -105
rect -497 -513 -463 -497
rect -401 -121 -367 -105
rect -401 -513 -367 -497
rect -305 -121 -271 -105
rect -305 -513 -271 -497
rect -209 -121 -175 -105
rect -209 -513 -175 -497
rect -113 -121 -79 -105
rect -113 -513 -79 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 79 -121 113 -105
rect 79 -513 113 -497
rect 175 -121 209 -105
rect 175 -513 209 -497
rect 271 -121 305 -105
rect 271 -513 305 -497
rect 367 -121 401 -105
rect 367 -513 401 -497
rect 463 -121 497 -105
rect 463 -513 497 -497
rect 559 -121 593 -105
rect 559 -513 593 -497
rect 655 -121 689 -105
rect 655 -513 689 -497
rect 751 -121 785 -105
rect 751 -513 785 -497
rect 847 -121 881 -105
rect 847 -513 881 -497
rect 943 -121 977 -105
rect 943 -513 977 -497
rect 1039 -121 1073 -105
rect 1039 -513 1073 -497
rect 1135 -121 1169 -105
rect 1135 -513 1169 -497
rect 1231 -121 1265 -105
rect 1231 -513 1265 -497
rect 1327 -121 1361 -105
rect 1327 -513 1361 -497
rect 1423 -121 1457 -105
rect 1423 -513 1457 -497
rect 1519 -121 1553 -105
rect 1519 -513 1553 -497
rect 1615 -121 1649 -105
rect 1615 -513 1649 -497
rect 1711 -121 1745 -105
rect 1711 -513 1745 -497
rect 1807 -121 1841 -105
rect 1807 -513 1841 -497
rect 1903 -121 1937 -105
rect 1903 -513 1937 -497
rect 1999 -121 2033 -105
rect 1999 -513 2033 -497
rect 2095 -121 2129 -105
rect 2095 -513 2129 -497
rect 2191 -121 2225 -105
rect 2191 -513 2225 -497
rect 2287 -121 2321 -105
rect 2287 -513 2321 -497
rect 2383 -121 2417 -105
rect 2383 -513 2417 -497
rect -2289 -581 -2273 -547
rect -2239 -581 -2223 -547
rect -2097 -581 -2081 -547
rect -2047 -581 -2031 -547
rect -1905 -581 -1889 -547
rect -1855 -581 -1839 -547
rect -1713 -581 -1697 -547
rect -1663 -581 -1647 -547
rect -1521 -581 -1505 -547
rect -1471 -581 -1455 -547
rect -1329 -581 -1313 -547
rect -1279 -581 -1263 -547
rect -1137 -581 -1121 -547
rect -1087 -581 -1071 -547
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 975 -581 991 -547
rect 1025 -581 1041 -547
rect 1167 -581 1183 -547
rect 1217 -581 1233 -547
rect 1359 -581 1375 -547
rect 1409 -581 1425 -547
rect 1551 -581 1567 -547
rect 1601 -581 1617 -547
rect 1743 -581 1759 -547
rect 1793 -581 1809 -547
rect 1935 -581 1951 -547
rect 1985 -581 2001 -547
rect 2127 -581 2143 -547
rect 2177 -581 2193 -547
rect 2319 -581 2335 -547
rect 2369 -581 2385 -547
rect -2289 -689 -2273 -655
rect -2239 -689 -2223 -655
rect -2097 -689 -2081 -655
rect -2047 -689 -2031 -655
rect -1905 -689 -1889 -655
rect -1855 -689 -1839 -655
rect -1713 -689 -1697 -655
rect -1663 -689 -1647 -655
rect -1521 -689 -1505 -655
rect -1471 -689 -1455 -655
rect -1329 -689 -1313 -655
rect -1279 -689 -1263 -655
rect -1137 -689 -1121 -655
rect -1087 -689 -1071 -655
rect -945 -689 -929 -655
rect -895 -689 -879 -655
rect -753 -689 -737 -655
rect -703 -689 -687 -655
rect -561 -689 -545 -655
rect -511 -689 -495 -655
rect -369 -689 -353 -655
rect -319 -689 -303 -655
rect -177 -689 -161 -655
rect -127 -689 -111 -655
rect 15 -689 31 -655
rect 65 -689 81 -655
rect 207 -689 223 -655
rect 257 -689 273 -655
rect 399 -689 415 -655
rect 449 -689 465 -655
rect 591 -689 607 -655
rect 641 -689 657 -655
rect 783 -689 799 -655
rect 833 -689 849 -655
rect 975 -689 991 -655
rect 1025 -689 1041 -655
rect 1167 -689 1183 -655
rect 1217 -689 1233 -655
rect 1359 -689 1375 -655
rect 1409 -689 1425 -655
rect 1551 -689 1567 -655
rect 1601 -689 1617 -655
rect 1743 -689 1759 -655
rect 1793 -689 1809 -655
rect 1935 -689 1951 -655
rect 1985 -689 2001 -655
rect 2127 -689 2143 -655
rect 2177 -689 2193 -655
rect 2319 -689 2335 -655
rect 2369 -689 2385 -655
rect -2417 -739 -2383 -723
rect -2417 -1131 -2383 -1115
rect -2321 -739 -2287 -723
rect -2321 -1131 -2287 -1115
rect -2225 -739 -2191 -723
rect -2225 -1131 -2191 -1115
rect -2129 -739 -2095 -723
rect -2129 -1131 -2095 -1115
rect -2033 -739 -1999 -723
rect -2033 -1131 -1999 -1115
rect -1937 -739 -1903 -723
rect -1937 -1131 -1903 -1115
rect -1841 -739 -1807 -723
rect -1841 -1131 -1807 -1115
rect -1745 -739 -1711 -723
rect -1745 -1131 -1711 -1115
rect -1649 -739 -1615 -723
rect -1649 -1131 -1615 -1115
rect -1553 -739 -1519 -723
rect -1553 -1131 -1519 -1115
rect -1457 -739 -1423 -723
rect -1457 -1131 -1423 -1115
rect -1361 -739 -1327 -723
rect -1361 -1131 -1327 -1115
rect -1265 -739 -1231 -723
rect -1265 -1131 -1231 -1115
rect -1169 -739 -1135 -723
rect -1169 -1131 -1135 -1115
rect -1073 -739 -1039 -723
rect -1073 -1131 -1039 -1115
rect -977 -739 -943 -723
rect -977 -1131 -943 -1115
rect -881 -739 -847 -723
rect -881 -1131 -847 -1115
rect -785 -739 -751 -723
rect -785 -1131 -751 -1115
rect -689 -739 -655 -723
rect -689 -1131 -655 -1115
rect -593 -739 -559 -723
rect -593 -1131 -559 -1115
rect -497 -739 -463 -723
rect -497 -1131 -463 -1115
rect -401 -739 -367 -723
rect -401 -1131 -367 -1115
rect -305 -739 -271 -723
rect -305 -1131 -271 -1115
rect -209 -739 -175 -723
rect -209 -1131 -175 -1115
rect -113 -739 -79 -723
rect -113 -1131 -79 -1115
rect -17 -739 17 -723
rect -17 -1131 17 -1115
rect 79 -739 113 -723
rect 79 -1131 113 -1115
rect 175 -739 209 -723
rect 175 -1131 209 -1115
rect 271 -739 305 -723
rect 271 -1131 305 -1115
rect 367 -739 401 -723
rect 367 -1131 401 -1115
rect 463 -739 497 -723
rect 463 -1131 497 -1115
rect 559 -739 593 -723
rect 559 -1131 593 -1115
rect 655 -739 689 -723
rect 655 -1131 689 -1115
rect 751 -739 785 -723
rect 751 -1131 785 -1115
rect 847 -739 881 -723
rect 847 -1131 881 -1115
rect 943 -739 977 -723
rect 943 -1131 977 -1115
rect 1039 -739 1073 -723
rect 1039 -1131 1073 -1115
rect 1135 -739 1169 -723
rect 1135 -1131 1169 -1115
rect 1231 -739 1265 -723
rect 1231 -1131 1265 -1115
rect 1327 -739 1361 -723
rect 1327 -1131 1361 -1115
rect 1423 -739 1457 -723
rect 1423 -1131 1457 -1115
rect 1519 -739 1553 -723
rect 1519 -1131 1553 -1115
rect 1615 -739 1649 -723
rect 1615 -1131 1649 -1115
rect 1711 -739 1745 -723
rect 1711 -1131 1745 -1115
rect 1807 -739 1841 -723
rect 1807 -1131 1841 -1115
rect 1903 -739 1937 -723
rect 1903 -1131 1937 -1115
rect 1999 -739 2033 -723
rect 1999 -1131 2033 -1115
rect 2095 -739 2129 -723
rect 2095 -1131 2129 -1115
rect 2191 -739 2225 -723
rect 2191 -1131 2225 -1115
rect 2287 -739 2321 -723
rect 2287 -1131 2321 -1115
rect 2383 -739 2417 -723
rect 2383 -1131 2417 -1115
rect -2385 -1199 -2369 -1165
rect -2335 -1199 -2319 -1165
rect -2193 -1199 -2177 -1165
rect -2143 -1199 -2127 -1165
rect -2001 -1199 -1985 -1165
rect -1951 -1199 -1935 -1165
rect -1809 -1199 -1793 -1165
rect -1759 -1199 -1743 -1165
rect -1617 -1199 -1601 -1165
rect -1567 -1199 -1551 -1165
rect -1425 -1199 -1409 -1165
rect -1375 -1199 -1359 -1165
rect -1233 -1199 -1217 -1165
rect -1183 -1199 -1167 -1165
rect -1041 -1199 -1025 -1165
rect -991 -1199 -975 -1165
rect -849 -1199 -833 -1165
rect -799 -1199 -783 -1165
rect -657 -1199 -641 -1165
rect -607 -1199 -591 -1165
rect -465 -1199 -449 -1165
rect -415 -1199 -399 -1165
rect -273 -1199 -257 -1165
rect -223 -1199 -207 -1165
rect -81 -1199 -65 -1165
rect -31 -1199 -15 -1165
rect 111 -1199 127 -1165
rect 161 -1199 177 -1165
rect 303 -1199 319 -1165
rect 353 -1199 369 -1165
rect 495 -1199 511 -1165
rect 545 -1199 561 -1165
rect 687 -1199 703 -1165
rect 737 -1199 753 -1165
rect 879 -1199 895 -1165
rect 929 -1199 945 -1165
rect 1071 -1199 1087 -1165
rect 1121 -1199 1137 -1165
rect 1263 -1199 1279 -1165
rect 1313 -1199 1329 -1165
rect 1455 -1199 1471 -1165
rect 1505 -1199 1521 -1165
rect 1647 -1199 1663 -1165
rect 1697 -1199 1713 -1165
rect 1839 -1199 1855 -1165
rect 1889 -1199 1905 -1165
rect 2031 -1199 2047 -1165
rect 2081 -1199 2097 -1165
rect 2223 -1199 2239 -1165
rect 2273 -1199 2289 -1165
rect -2531 -1267 -2497 -1205
rect 2497 -1267 2531 -1205
rect -2531 -1301 -2435 -1267
rect 2435 -1301 2531 -1267
<< viali >>
rect -2369 1165 -2335 1199
rect -2177 1165 -2143 1199
rect -1985 1165 -1951 1199
rect -1793 1165 -1759 1199
rect -1601 1165 -1567 1199
rect -1409 1165 -1375 1199
rect -1217 1165 -1183 1199
rect -1025 1165 -991 1199
rect -833 1165 -799 1199
rect -641 1165 -607 1199
rect -449 1165 -415 1199
rect -257 1165 -223 1199
rect -65 1165 -31 1199
rect 127 1165 161 1199
rect 319 1165 353 1199
rect 511 1165 545 1199
rect 703 1165 737 1199
rect 895 1165 929 1199
rect 1087 1165 1121 1199
rect 1279 1165 1313 1199
rect 1471 1165 1505 1199
rect 1663 1165 1697 1199
rect 1855 1165 1889 1199
rect 2047 1165 2081 1199
rect 2239 1165 2273 1199
rect -2417 739 -2383 1115
rect -2321 739 -2287 1115
rect -2225 739 -2191 1115
rect -2129 739 -2095 1115
rect -2033 739 -1999 1115
rect -1937 739 -1903 1115
rect -1841 739 -1807 1115
rect -1745 739 -1711 1115
rect -1649 739 -1615 1115
rect -1553 739 -1519 1115
rect -1457 739 -1423 1115
rect -1361 739 -1327 1115
rect -1265 739 -1231 1115
rect -1169 739 -1135 1115
rect -1073 739 -1039 1115
rect -977 739 -943 1115
rect -881 739 -847 1115
rect -785 739 -751 1115
rect -689 739 -655 1115
rect -593 739 -559 1115
rect -497 739 -463 1115
rect -401 739 -367 1115
rect -305 739 -271 1115
rect -209 739 -175 1115
rect -113 739 -79 1115
rect -17 739 17 1115
rect 79 739 113 1115
rect 175 739 209 1115
rect 271 739 305 1115
rect 367 739 401 1115
rect 463 739 497 1115
rect 559 739 593 1115
rect 655 739 689 1115
rect 751 739 785 1115
rect 847 739 881 1115
rect 943 739 977 1115
rect 1039 739 1073 1115
rect 1135 739 1169 1115
rect 1231 739 1265 1115
rect 1327 739 1361 1115
rect 1423 739 1457 1115
rect 1519 739 1553 1115
rect 1615 739 1649 1115
rect 1711 739 1745 1115
rect 1807 739 1841 1115
rect 1903 739 1937 1115
rect 1999 739 2033 1115
rect 2095 739 2129 1115
rect 2191 739 2225 1115
rect 2287 739 2321 1115
rect 2383 739 2417 1115
rect -2273 655 -2239 689
rect -2081 655 -2047 689
rect -1889 655 -1855 689
rect -1697 655 -1663 689
rect -1505 655 -1471 689
rect -1313 655 -1279 689
rect -1121 655 -1087 689
rect -929 655 -895 689
rect -737 655 -703 689
rect -545 655 -511 689
rect -353 655 -319 689
rect -161 655 -127 689
rect 31 655 65 689
rect 223 655 257 689
rect 415 655 449 689
rect 607 655 641 689
rect 799 655 833 689
rect 991 655 1025 689
rect 1183 655 1217 689
rect 1375 655 1409 689
rect 1567 655 1601 689
rect 1759 655 1793 689
rect 1951 655 1985 689
rect 2143 655 2177 689
rect 2335 655 2369 689
rect -2273 547 -2239 581
rect -2081 547 -2047 581
rect -1889 547 -1855 581
rect -1697 547 -1663 581
rect -1505 547 -1471 581
rect -1313 547 -1279 581
rect -1121 547 -1087 581
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect 991 547 1025 581
rect 1183 547 1217 581
rect 1375 547 1409 581
rect 1567 547 1601 581
rect 1759 547 1793 581
rect 1951 547 1985 581
rect 2143 547 2177 581
rect 2335 547 2369 581
rect -2417 121 -2383 497
rect -2321 121 -2287 497
rect -2225 121 -2191 497
rect -2129 121 -2095 497
rect -2033 121 -1999 497
rect -1937 121 -1903 497
rect -1841 121 -1807 497
rect -1745 121 -1711 497
rect -1649 121 -1615 497
rect -1553 121 -1519 497
rect -1457 121 -1423 497
rect -1361 121 -1327 497
rect -1265 121 -1231 497
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect 1231 121 1265 497
rect 1327 121 1361 497
rect 1423 121 1457 497
rect 1519 121 1553 497
rect 1615 121 1649 497
rect 1711 121 1745 497
rect 1807 121 1841 497
rect 1903 121 1937 497
rect 1999 121 2033 497
rect 2095 121 2129 497
rect 2191 121 2225 497
rect 2287 121 2321 497
rect 2383 121 2417 497
rect -2369 37 -2335 71
rect -2177 37 -2143 71
rect -1985 37 -1951 71
rect -1793 37 -1759 71
rect -1601 37 -1567 71
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect 1471 37 1505 71
rect 1663 37 1697 71
rect 1855 37 1889 71
rect 2047 37 2081 71
rect 2239 37 2273 71
rect -2369 -71 -2335 -37
rect -2177 -71 -2143 -37
rect -1985 -71 -1951 -37
rect -1793 -71 -1759 -37
rect -1601 -71 -1567 -37
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect 1471 -71 1505 -37
rect 1663 -71 1697 -37
rect 1855 -71 1889 -37
rect 2047 -71 2081 -37
rect 2239 -71 2273 -37
rect -2417 -497 -2383 -121
rect -2321 -497 -2287 -121
rect -2225 -497 -2191 -121
rect -2129 -497 -2095 -121
rect -2033 -497 -1999 -121
rect -1937 -497 -1903 -121
rect -1841 -497 -1807 -121
rect -1745 -497 -1711 -121
rect -1649 -497 -1615 -121
rect -1553 -497 -1519 -121
rect -1457 -497 -1423 -121
rect -1361 -497 -1327 -121
rect -1265 -497 -1231 -121
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect 1231 -497 1265 -121
rect 1327 -497 1361 -121
rect 1423 -497 1457 -121
rect 1519 -497 1553 -121
rect 1615 -497 1649 -121
rect 1711 -497 1745 -121
rect 1807 -497 1841 -121
rect 1903 -497 1937 -121
rect 1999 -497 2033 -121
rect 2095 -497 2129 -121
rect 2191 -497 2225 -121
rect 2287 -497 2321 -121
rect 2383 -497 2417 -121
rect -2273 -581 -2239 -547
rect -2081 -581 -2047 -547
rect -1889 -581 -1855 -547
rect -1697 -581 -1663 -547
rect -1505 -581 -1471 -547
rect -1313 -581 -1279 -547
rect -1121 -581 -1087 -547
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
rect 991 -581 1025 -547
rect 1183 -581 1217 -547
rect 1375 -581 1409 -547
rect 1567 -581 1601 -547
rect 1759 -581 1793 -547
rect 1951 -581 1985 -547
rect 2143 -581 2177 -547
rect 2335 -581 2369 -547
rect -2273 -689 -2239 -655
rect -2081 -689 -2047 -655
rect -1889 -689 -1855 -655
rect -1697 -689 -1663 -655
rect -1505 -689 -1471 -655
rect -1313 -689 -1279 -655
rect -1121 -689 -1087 -655
rect -929 -689 -895 -655
rect -737 -689 -703 -655
rect -545 -689 -511 -655
rect -353 -689 -319 -655
rect -161 -689 -127 -655
rect 31 -689 65 -655
rect 223 -689 257 -655
rect 415 -689 449 -655
rect 607 -689 641 -655
rect 799 -689 833 -655
rect 991 -689 1025 -655
rect 1183 -689 1217 -655
rect 1375 -689 1409 -655
rect 1567 -689 1601 -655
rect 1759 -689 1793 -655
rect 1951 -689 1985 -655
rect 2143 -689 2177 -655
rect 2335 -689 2369 -655
rect -2417 -1115 -2383 -739
rect -2321 -1115 -2287 -739
rect -2225 -1115 -2191 -739
rect -2129 -1115 -2095 -739
rect -2033 -1115 -1999 -739
rect -1937 -1115 -1903 -739
rect -1841 -1115 -1807 -739
rect -1745 -1115 -1711 -739
rect -1649 -1115 -1615 -739
rect -1553 -1115 -1519 -739
rect -1457 -1115 -1423 -739
rect -1361 -1115 -1327 -739
rect -1265 -1115 -1231 -739
rect -1169 -1115 -1135 -739
rect -1073 -1115 -1039 -739
rect -977 -1115 -943 -739
rect -881 -1115 -847 -739
rect -785 -1115 -751 -739
rect -689 -1115 -655 -739
rect -593 -1115 -559 -739
rect -497 -1115 -463 -739
rect -401 -1115 -367 -739
rect -305 -1115 -271 -739
rect -209 -1115 -175 -739
rect -113 -1115 -79 -739
rect -17 -1115 17 -739
rect 79 -1115 113 -739
rect 175 -1115 209 -739
rect 271 -1115 305 -739
rect 367 -1115 401 -739
rect 463 -1115 497 -739
rect 559 -1115 593 -739
rect 655 -1115 689 -739
rect 751 -1115 785 -739
rect 847 -1115 881 -739
rect 943 -1115 977 -739
rect 1039 -1115 1073 -739
rect 1135 -1115 1169 -739
rect 1231 -1115 1265 -739
rect 1327 -1115 1361 -739
rect 1423 -1115 1457 -739
rect 1519 -1115 1553 -739
rect 1615 -1115 1649 -739
rect 1711 -1115 1745 -739
rect 1807 -1115 1841 -739
rect 1903 -1115 1937 -739
rect 1999 -1115 2033 -739
rect 2095 -1115 2129 -739
rect 2191 -1115 2225 -739
rect 2287 -1115 2321 -739
rect 2383 -1115 2417 -739
rect -2369 -1199 -2335 -1165
rect -2177 -1199 -2143 -1165
rect -1985 -1199 -1951 -1165
rect -1793 -1199 -1759 -1165
rect -1601 -1199 -1567 -1165
rect -1409 -1199 -1375 -1165
rect -1217 -1199 -1183 -1165
rect -1025 -1199 -991 -1165
rect -833 -1199 -799 -1165
rect -641 -1199 -607 -1165
rect -449 -1199 -415 -1165
rect -257 -1199 -223 -1165
rect -65 -1199 -31 -1165
rect 127 -1199 161 -1165
rect 319 -1199 353 -1165
rect 511 -1199 545 -1165
rect 703 -1199 737 -1165
rect 895 -1199 929 -1165
rect 1087 -1199 1121 -1165
rect 1279 -1199 1313 -1165
rect 1471 -1199 1505 -1165
rect 1663 -1199 1697 -1165
rect 1855 -1199 1889 -1165
rect 2047 -1199 2081 -1165
rect 2239 -1199 2273 -1165
<< metal1 >>
rect -2381 1199 -2323 1205
rect -2381 1165 -2369 1199
rect -2335 1165 -2323 1199
rect -2381 1159 -2323 1165
rect -2189 1199 -2131 1205
rect -2189 1165 -2177 1199
rect -2143 1165 -2131 1199
rect -2189 1159 -2131 1165
rect -1997 1199 -1939 1205
rect -1997 1165 -1985 1199
rect -1951 1165 -1939 1199
rect -1997 1159 -1939 1165
rect -1805 1199 -1747 1205
rect -1805 1165 -1793 1199
rect -1759 1165 -1747 1199
rect -1805 1159 -1747 1165
rect -1613 1199 -1555 1205
rect -1613 1165 -1601 1199
rect -1567 1165 -1555 1199
rect -1613 1159 -1555 1165
rect -1421 1199 -1363 1205
rect -1421 1165 -1409 1199
rect -1375 1165 -1363 1199
rect -1421 1159 -1363 1165
rect -1229 1199 -1171 1205
rect -1229 1165 -1217 1199
rect -1183 1165 -1171 1199
rect -1229 1159 -1171 1165
rect -1037 1199 -979 1205
rect -1037 1165 -1025 1199
rect -991 1165 -979 1199
rect -1037 1159 -979 1165
rect -845 1199 -787 1205
rect -845 1165 -833 1199
rect -799 1165 -787 1199
rect -845 1159 -787 1165
rect -653 1199 -595 1205
rect -653 1165 -641 1199
rect -607 1165 -595 1199
rect -653 1159 -595 1165
rect -461 1199 -403 1205
rect -461 1165 -449 1199
rect -415 1165 -403 1199
rect -461 1159 -403 1165
rect -269 1199 -211 1205
rect -269 1165 -257 1199
rect -223 1165 -211 1199
rect -269 1159 -211 1165
rect -77 1199 -19 1205
rect -77 1165 -65 1199
rect -31 1165 -19 1199
rect -77 1159 -19 1165
rect 115 1199 173 1205
rect 115 1165 127 1199
rect 161 1165 173 1199
rect 115 1159 173 1165
rect 307 1199 365 1205
rect 307 1165 319 1199
rect 353 1165 365 1199
rect 307 1159 365 1165
rect 499 1199 557 1205
rect 499 1165 511 1199
rect 545 1165 557 1199
rect 499 1159 557 1165
rect 691 1199 749 1205
rect 691 1165 703 1199
rect 737 1165 749 1199
rect 691 1159 749 1165
rect 883 1199 941 1205
rect 883 1165 895 1199
rect 929 1165 941 1199
rect 883 1159 941 1165
rect 1075 1199 1133 1205
rect 1075 1165 1087 1199
rect 1121 1165 1133 1199
rect 1075 1159 1133 1165
rect 1267 1199 1325 1205
rect 1267 1165 1279 1199
rect 1313 1165 1325 1199
rect 1267 1159 1325 1165
rect 1459 1199 1517 1205
rect 1459 1165 1471 1199
rect 1505 1165 1517 1199
rect 1459 1159 1517 1165
rect 1651 1199 1709 1205
rect 1651 1165 1663 1199
rect 1697 1165 1709 1199
rect 1651 1159 1709 1165
rect 1843 1199 1901 1205
rect 1843 1165 1855 1199
rect 1889 1165 1901 1199
rect 1843 1159 1901 1165
rect 2035 1199 2093 1205
rect 2035 1165 2047 1199
rect 2081 1165 2093 1199
rect 2035 1159 2093 1165
rect 2227 1199 2285 1205
rect 2227 1165 2239 1199
rect 2273 1165 2285 1199
rect 2227 1159 2285 1165
rect -2423 1115 -2377 1127
rect -2423 739 -2417 1115
rect -2383 739 -2377 1115
rect -2423 727 -2377 739
rect -2327 1115 -2281 1127
rect -2327 739 -2321 1115
rect -2287 739 -2281 1115
rect -2327 727 -2281 739
rect -2231 1115 -2185 1127
rect -2231 739 -2225 1115
rect -2191 739 -2185 1115
rect -2231 727 -2185 739
rect -2135 1115 -2089 1127
rect -2135 739 -2129 1115
rect -2095 739 -2089 1115
rect -2135 727 -2089 739
rect -2039 1115 -1993 1127
rect -2039 739 -2033 1115
rect -1999 739 -1993 1115
rect -2039 727 -1993 739
rect -1943 1115 -1897 1127
rect -1943 739 -1937 1115
rect -1903 739 -1897 1115
rect -1943 727 -1897 739
rect -1847 1115 -1801 1127
rect -1847 739 -1841 1115
rect -1807 739 -1801 1115
rect -1847 727 -1801 739
rect -1751 1115 -1705 1127
rect -1751 739 -1745 1115
rect -1711 739 -1705 1115
rect -1751 727 -1705 739
rect -1655 1115 -1609 1127
rect -1655 739 -1649 1115
rect -1615 739 -1609 1115
rect -1655 727 -1609 739
rect -1559 1115 -1513 1127
rect -1559 739 -1553 1115
rect -1519 739 -1513 1115
rect -1559 727 -1513 739
rect -1463 1115 -1417 1127
rect -1463 739 -1457 1115
rect -1423 739 -1417 1115
rect -1463 727 -1417 739
rect -1367 1115 -1321 1127
rect -1367 739 -1361 1115
rect -1327 739 -1321 1115
rect -1367 727 -1321 739
rect -1271 1115 -1225 1127
rect -1271 739 -1265 1115
rect -1231 739 -1225 1115
rect -1271 727 -1225 739
rect -1175 1115 -1129 1127
rect -1175 739 -1169 1115
rect -1135 739 -1129 1115
rect -1175 727 -1129 739
rect -1079 1115 -1033 1127
rect -1079 739 -1073 1115
rect -1039 739 -1033 1115
rect -1079 727 -1033 739
rect -983 1115 -937 1127
rect -983 739 -977 1115
rect -943 739 -937 1115
rect -983 727 -937 739
rect -887 1115 -841 1127
rect -887 739 -881 1115
rect -847 739 -841 1115
rect -887 727 -841 739
rect -791 1115 -745 1127
rect -791 739 -785 1115
rect -751 739 -745 1115
rect -791 727 -745 739
rect -695 1115 -649 1127
rect -695 739 -689 1115
rect -655 739 -649 1115
rect -695 727 -649 739
rect -599 1115 -553 1127
rect -599 739 -593 1115
rect -559 739 -553 1115
rect -599 727 -553 739
rect -503 1115 -457 1127
rect -503 739 -497 1115
rect -463 739 -457 1115
rect -503 727 -457 739
rect -407 1115 -361 1127
rect -407 739 -401 1115
rect -367 739 -361 1115
rect -407 727 -361 739
rect -311 1115 -265 1127
rect -311 739 -305 1115
rect -271 739 -265 1115
rect -311 727 -265 739
rect -215 1115 -169 1127
rect -215 739 -209 1115
rect -175 739 -169 1115
rect -215 727 -169 739
rect -119 1115 -73 1127
rect -119 739 -113 1115
rect -79 739 -73 1115
rect -119 727 -73 739
rect -23 1115 23 1127
rect -23 739 -17 1115
rect 17 739 23 1115
rect -23 727 23 739
rect 73 1115 119 1127
rect 73 739 79 1115
rect 113 739 119 1115
rect 73 727 119 739
rect 169 1115 215 1127
rect 169 739 175 1115
rect 209 739 215 1115
rect 169 727 215 739
rect 265 1115 311 1127
rect 265 739 271 1115
rect 305 739 311 1115
rect 265 727 311 739
rect 361 1115 407 1127
rect 361 739 367 1115
rect 401 739 407 1115
rect 361 727 407 739
rect 457 1115 503 1127
rect 457 739 463 1115
rect 497 739 503 1115
rect 457 727 503 739
rect 553 1115 599 1127
rect 553 739 559 1115
rect 593 739 599 1115
rect 553 727 599 739
rect 649 1115 695 1127
rect 649 739 655 1115
rect 689 739 695 1115
rect 649 727 695 739
rect 745 1115 791 1127
rect 745 739 751 1115
rect 785 739 791 1115
rect 745 727 791 739
rect 841 1115 887 1127
rect 841 739 847 1115
rect 881 739 887 1115
rect 841 727 887 739
rect 937 1115 983 1127
rect 937 739 943 1115
rect 977 739 983 1115
rect 937 727 983 739
rect 1033 1115 1079 1127
rect 1033 739 1039 1115
rect 1073 739 1079 1115
rect 1033 727 1079 739
rect 1129 1115 1175 1127
rect 1129 739 1135 1115
rect 1169 739 1175 1115
rect 1129 727 1175 739
rect 1225 1115 1271 1127
rect 1225 739 1231 1115
rect 1265 739 1271 1115
rect 1225 727 1271 739
rect 1321 1115 1367 1127
rect 1321 739 1327 1115
rect 1361 739 1367 1115
rect 1321 727 1367 739
rect 1417 1115 1463 1127
rect 1417 739 1423 1115
rect 1457 739 1463 1115
rect 1417 727 1463 739
rect 1513 1115 1559 1127
rect 1513 739 1519 1115
rect 1553 739 1559 1115
rect 1513 727 1559 739
rect 1609 1115 1655 1127
rect 1609 739 1615 1115
rect 1649 739 1655 1115
rect 1609 727 1655 739
rect 1705 1115 1751 1127
rect 1705 739 1711 1115
rect 1745 739 1751 1115
rect 1705 727 1751 739
rect 1801 1115 1847 1127
rect 1801 739 1807 1115
rect 1841 739 1847 1115
rect 1801 727 1847 739
rect 1897 1115 1943 1127
rect 1897 739 1903 1115
rect 1937 739 1943 1115
rect 1897 727 1943 739
rect 1993 1115 2039 1127
rect 1993 739 1999 1115
rect 2033 739 2039 1115
rect 1993 727 2039 739
rect 2089 1115 2135 1127
rect 2089 739 2095 1115
rect 2129 739 2135 1115
rect 2089 727 2135 739
rect 2185 1115 2231 1127
rect 2185 739 2191 1115
rect 2225 739 2231 1115
rect 2185 727 2231 739
rect 2281 1115 2327 1127
rect 2281 739 2287 1115
rect 2321 739 2327 1115
rect 2281 727 2327 739
rect 2377 1115 2423 1127
rect 2377 739 2383 1115
rect 2417 739 2423 1115
rect 2377 727 2423 739
rect -2285 689 -2227 695
rect -2285 655 -2273 689
rect -2239 655 -2227 689
rect -2285 649 -2227 655
rect -2093 689 -2035 695
rect -2093 655 -2081 689
rect -2047 655 -2035 689
rect -2093 649 -2035 655
rect -1901 689 -1843 695
rect -1901 655 -1889 689
rect -1855 655 -1843 689
rect -1901 649 -1843 655
rect -1709 689 -1651 695
rect -1709 655 -1697 689
rect -1663 655 -1651 689
rect -1709 649 -1651 655
rect -1517 689 -1459 695
rect -1517 655 -1505 689
rect -1471 655 -1459 689
rect -1517 649 -1459 655
rect -1325 689 -1267 695
rect -1325 655 -1313 689
rect -1279 655 -1267 689
rect -1325 649 -1267 655
rect -1133 689 -1075 695
rect -1133 655 -1121 689
rect -1087 655 -1075 689
rect -1133 649 -1075 655
rect -941 689 -883 695
rect -941 655 -929 689
rect -895 655 -883 689
rect -941 649 -883 655
rect -749 689 -691 695
rect -749 655 -737 689
rect -703 655 -691 689
rect -749 649 -691 655
rect -557 689 -499 695
rect -557 655 -545 689
rect -511 655 -499 689
rect -557 649 -499 655
rect -365 689 -307 695
rect -365 655 -353 689
rect -319 655 -307 689
rect -365 649 -307 655
rect -173 689 -115 695
rect -173 655 -161 689
rect -127 655 -115 689
rect -173 649 -115 655
rect 19 689 77 695
rect 19 655 31 689
rect 65 655 77 689
rect 19 649 77 655
rect 211 689 269 695
rect 211 655 223 689
rect 257 655 269 689
rect 211 649 269 655
rect 403 689 461 695
rect 403 655 415 689
rect 449 655 461 689
rect 403 649 461 655
rect 595 689 653 695
rect 595 655 607 689
rect 641 655 653 689
rect 595 649 653 655
rect 787 689 845 695
rect 787 655 799 689
rect 833 655 845 689
rect 787 649 845 655
rect 979 689 1037 695
rect 979 655 991 689
rect 1025 655 1037 689
rect 979 649 1037 655
rect 1171 689 1229 695
rect 1171 655 1183 689
rect 1217 655 1229 689
rect 1171 649 1229 655
rect 1363 689 1421 695
rect 1363 655 1375 689
rect 1409 655 1421 689
rect 1363 649 1421 655
rect 1555 689 1613 695
rect 1555 655 1567 689
rect 1601 655 1613 689
rect 1555 649 1613 655
rect 1747 689 1805 695
rect 1747 655 1759 689
rect 1793 655 1805 689
rect 1747 649 1805 655
rect 1939 689 1997 695
rect 1939 655 1951 689
rect 1985 655 1997 689
rect 1939 649 1997 655
rect 2131 689 2189 695
rect 2131 655 2143 689
rect 2177 655 2189 689
rect 2131 649 2189 655
rect 2323 689 2381 695
rect 2323 655 2335 689
rect 2369 655 2381 689
rect 2323 649 2381 655
rect -2285 581 -2227 587
rect -2285 547 -2273 581
rect -2239 547 -2227 581
rect -2285 541 -2227 547
rect -2093 581 -2035 587
rect -2093 547 -2081 581
rect -2047 547 -2035 581
rect -2093 541 -2035 547
rect -1901 581 -1843 587
rect -1901 547 -1889 581
rect -1855 547 -1843 581
rect -1901 541 -1843 547
rect -1709 581 -1651 587
rect -1709 547 -1697 581
rect -1663 547 -1651 581
rect -1709 541 -1651 547
rect -1517 581 -1459 587
rect -1517 547 -1505 581
rect -1471 547 -1459 581
rect -1517 541 -1459 547
rect -1325 581 -1267 587
rect -1325 547 -1313 581
rect -1279 547 -1267 581
rect -1325 541 -1267 547
rect -1133 581 -1075 587
rect -1133 547 -1121 581
rect -1087 547 -1075 581
rect -1133 541 -1075 547
rect -941 581 -883 587
rect -941 547 -929 581
rect -895 547 -883 581
rect -941 541 -883 547
rect -749 581 -691 587
rect -749 547 -737 581
rect -703 547 -691 581
rect -749 541 -691 547
rect -557 581 -499 587
rect -557 547 -545 581
rect -511 547 -499 581
rect -557 541 -499 547
rect -365 581 -307 587
rect -365 547 -353 581
rect -319 547 -307 581
rect -365 541 -307 547
rect -173 581 -115 587
rect -173 547 -161 581
rect -127 547 -115 581
rect -173 541 -115 547
rect 19 581 77 587
rect 19 547 31 581
rect 65 547 77 581
rect 19 541 77 547
rect 211 581 269 587
rect 211 547 223 581
rect 257 547 269 581
rect 211 541 269 547
rect 403 581 461 587
rect 403 547 415 581
rect 449 547 461 581
rect 403 541 461 547
rect 595 581 653 587
rect 595 547 607 581
rect 641 547 653 581
rect 595 541 653 547
rect 787 581 845 587
rect 787 547 799 581
rect 833 547 845 581
rect 787 541 845 547
rect 979 581 1037 587
rect 979 547 991 581
rect 1025 547 1037 581
rect 979 541 1037 547
rect 1171 581 1229 587
rect 1171 547 1183 581
rect 1217 547 1229 581
rect 1171 541 1229 547
rect 1363 581 1421 587
rect 1363 547 1375 581
rect 1409 547 1421 581
rect 1363 541 1421 547
rect 1555 581 1613 587
rect 1555 547 1567 581
rect 1601 547 1613 581
rect 1555 541 1613 547
rect 1747 581 1805 587
rect 1747 547 1759 581
rect 1793 547 1805 581
rect 1747 541 1805 547
rect 1939 581 1997 587
rect 1939 547 1951 581
rect 1985 547 1997 581
rect 1939 541 1997 547
rect 2131 581 2189 587
rect 2131 547 2143 581
rect 2177 547 2189 581
rect 2131 541 2189 547
rect 2323 581 2381 587
rect 2323 547 2335 581
rect 2369 547 2381 581
rect 2323 541 2381 547
rect -2423 497 -2377 509
rect -2423 121 -2417 497
rect -2383 121 -2377 497
rect -2423 109 -2377 121
rect -2327 497 -2281 509
rect -2327 121 -2321 497
rect -2287 121 -2281 497
rect -2327 109 -2281 121
rect -2231 497 -2185 509
rect -2231 121 -2225 497
rect -2191 121 -2185 497
rect -2231 109 -2185 121
rect -2135 497 -2089 509
rect -2135 121 -2129 497
rect -2095 121 -2089 497
rect -2135 109 -2089 121
rect -2039 497 -1993 509
rect -2039 121 -2033 497
rect -1999 121 -1993 497
rect -2039 109 -1993 121
rect -1943 497 -1897 509
rect -1943 121 -1937 497
rect -1903 121 -1897 497
rect -1943 109 -1897 121
rect -1847 497 -1801 509
rect -1847 121 -1841 497
rect -1807 121 -1801 497
rect -1847 109 -1801 121
rect -1751 497 -1705 509
rect -1751 121 -1745 497
rect -1711 121 -1705 497
rect -1751 109 -1705 121
rect -1655 497 -1609 509
rect -1655 121 -1649 497
rect -1615 121 -1609 497
rect -1655 109 -1609 121
rect -1559 497 -1513 509
rect -1559 121 -1553 497
rect -1519 121 -1513 497
rect -1559 109 -1513 121
rect -1463 497 -1417 509
rect -1463 121 -1457 497
rect -1423 121 -1417 497
rect -1463 109 -1417 121
rect -1367 497 -1321 509
rect -1367 121 -1361 497
rect -1327 121 -1321 497
rect -1367 109 -1321 121
rect -1271 497 -1225 509
rect -1271 121 -1265 497
rect -1231 121 -1225 497
rect -1271 109 -1225 121
rect -1175 497 -1129 509
rect -1175 121 -1169 497
rect -1135 121 -1129 497
rect -1175 109 -1129 121
rect -1079 497 -1033 509
rect -1079 121 -1073 497
rect -1039 121 -1033 497
rect -1079 109 -1033 121
rect -983 497 -937 509
rect -983 121 -977 497
rect -943 121 -937 497
rect -983 109 -937 121
rect -887 497 -841 509
rect -887 121 -881 497
rect -847 121 -841 497
rect -887 109 -841 121
rect -791 497 -745 509
rect -791 121 -785 497
rect -751 121 -745 497
rect -791 109 -745 121
rect -695 497 -649 509
rect -695 121 -689 497
rect -655 121 -649 497
rect -695 109 -649 121
rect -599 497 -553 509
rect -599 121 -593 497
rect -559 121 -553 497
rect -599 109 -553 121
rect -503 497 -457 509
rect -503 121 -497 497
rect -463 121 -457 497
rect -503 109 -457 121
rect -407 497 -361 509
rect -407 121 -401 497
rect -367 121 -361 497
rect -407 109 -361 121
rect -311 497 -265 509
rect -311 121 -305 497
rect -271 121 -265 497
rect -311 109 -265 121
rect -215 497 -169 509
rect -215 121 -209 497
rect -175 121 -169 497
rect -215 109 -169 121
rect -119 497 -73 509
rect -119 121 -113 497
rect -79 121 -73 497
rect -119 109 -73 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 73 497 119 509
rect 73 121 79 497
rect 113 121 119 497
rect 73 109 119 121
rect 169 497 215 509
rect 169 121 175 497
rect 209 121 215 497
rect 169 109 215 121
rect 265 497 311 509
rect 265 121 271 497
rect 305 121 311 497
rect 265 109 311 121
rect 361 497 407 509
rect 361 121 367 497
rect 401 121 407 497
rect 361 109 407 121
rect 457 497 503 509
rect 457 121 463 497
rect 497 121 503 497
rect 457 109 503 121
rect 553 497 599 509
rect 553 121 559 497
rect 593 121 599 497
rect 553 109 599 121
rect 649 497 695 509
rect 649 121 655 497
rect 689 121 695 497
rect 649 109 695 121
rect 745 497 791 509
rect 745 121 751 497
rect 785 121 791 497
rect 745 109 791 121
rect 841 497 887 509
rect 841 121 847 497
rect 881 121 887 497
rect 841 109 887 121
rect 937 497 983 509
rect 937 121 943 497
rect 977 121 983 497
rect 937 109 983 121
rect 1033 497 1079 509
rect 1033 121 1039 497
rect 1073 121 1079 497
rect 1033 109 1079 121
rect 1129 497 1175 509
rect 1129 121 1135 497
rect 1169 121 1175 497
rect 1129 109 1175 121
rect 1225 497 1271 509
rect 1225 121 1231 497
rect 1265 121 1271 497
rect 1225 109 1271 121
rect 1321 497 1367 509
rect 1321 121 1327 497
rect 1361 121 1367 497
rect 1321 109 1367 121
rect 1417 497 1463 509
rect 1417 121 1423 497
rect 1457 121 1463 497
rect 1417 109 1463 121
rect 1513 497 1559 509
rect 1513 121 1519 497
rect 1553 121 1559 497
rect 1513 109 1559 121
rect 1609 497 1655 509
rect 1609 121 1615 497
rect 1649 121 1655 497
rect 1609 109 1655 121
rect 1705 497 1751 509
rect 1705 121 1711 497
rect 1745 121 1751 497
rect 1705 109 1751 121
rect 1801 497 1847 509
rect 1801 121 1807 497
rect 1841 121 1847 497
rect 1801 109 1847 121
rect 1897 497 1943 509
rect 1897 121 1903 497
rect 1937 121 1943 497
rect 1897 109 1943 121
rect 1993 497 2039 509
rect 1993 121 1999 497
rect 2033 121 2039 497
rect 1993 109 2039 121
rect 2089 497 2135 509
rect 2089 121 2095 497
rect 2129 121 2135 497
rect 2089 109 2135 121
rect 2185 497 2231 509
rect 2185 121 2191 497
rect 2225 121 2231 497
rect 2185 109 2231 121
rect 2281 497 2327 509
rect 2281 121 2287 497
rect 2321 121 2327 497
rect 2281 109 2327 121
rect 2377 497 2423 509
rect 2377 121 2383 497
rect 2417 121 2423 497
rect 2377 109 2423 121
rect -2381 71 -2323 77
rect -2381 37 -2369 71
rect -2335 37 -2323 71
rect -2381 31 -2323 37
rect -2189 71 -2131 77
rect -2189 37 -2177 71
rect -2143 37 -2131 71
rect -2189 31 -2131 37
rect -1997 71 -1939 77
rect -1997 37 -1985 71
rect -1951 37 -1939 71
rect -1997 31 -1939 37
rect -1805 71 -1747 77
rect -1805 37 -1793 71
rect -1759 37 -1747 71
rect -1805 31 -1747 37
rect -1613 71 -1555 77
rect -1613 37 -1601 71
rect -1567 37 -1555 71
rect -1613 31 -1555 37
rect -1421 71 -1363 77
rect -1421 37 -1409 71
rect -1375 37 -1363 71
rect -1421 31 -1363 37
rect -1229 71 -1171 77
rect -1229 37 -1217 71
rect -1183 37 -1171 71
rect -1229 31 -1171 37
rect -1037 71 -979 77
rect -1037 37 -1025 71
rect -991 37 -979 71
rect -1037 31 -979 37
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect 1075 71 1133 77
rect 1075 37 1087 71
rect 1121 37 1133 71
rect 1075 31 1133 37
rect 1267 71 1325 77
rect 1267 37 1279 71
rect 1313 37 1325 71
rect 1267 31 1325 37
rect 1459 71 1517 77
rect 1459 37 1471 71
rect 1505 37 1517 71
rect 1459 31 1517 37
rect 1651 71 1709 77
rect 1651 37 1663 71
rect 1697 37 1709 71
rect 1651 31 1709 37
rect 1843 71 1901 77
rect 1843 37 1855 71
rect 1889 37 1901 71
rect 1843 31 1901 37
rect 2035 71 2093 77
rect 2035 37 2047 71
rect 2081 37 2093 71
rect 2035 31 2093 37
rect 2227 71 2285 77
rect 2227 37 2239 71
rect 2273 37 2285 71
rect 2227 31 2285 37
rect -2381 -37 -2323 -31
rect -2381 -71 -2369 -37
rect -2335 -71 -2323 -37
rect -2381 -77 -2323 -71
rect -2189 -37 -2131 -31
rect -2189 -71 -2177 -37
rect -2143 -71 -2131 -37
rect -2189 -77 -2131 -71
rect -1997 -37 -1939 -31
rect -1997 -71 -1985 -37
rect -1951 -71 -1939 -37
rect -1997 -77 -1939 -71
rect -1805 -37 -1747 -31
rect -1805 -71 -1793 -37
rect -1759 -71 -1747 -37
rect -1805 -77 -1747 -71
rect -1613 -37 -1555 -31
rect -1613 -71 -1601 -37
rect -1567 -71 -1555 -37
rect -1613 -77 -1555 -71
rect -1421 -37 -1363 -31
rect -1421 -71 -1409 -37
rect -1375 -71 -1363 -37
rect -1421 -77 -1363 -71
rect -1229 -37 -1171 -31
rect -1229 -71 -1217 -37
rect -1183 -71 -1171 -37
rect -1229 -77 -1171 -71
rect -1037 -37 -979 -31
rect -1037 -71 -1025 -37
rect -991 -71 -979 -37
rect -1037 -77 -979 -71
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect 1075 -37 1133 -31
rect 1075 -71 1087 -37
rect 1121 -71 1133 -37
rect 1075 -77 1133 -71
rect 1267 -37 1325 -31
rect 1267 -71 1279 -37
rect 1313 -71 1325 -37
rect 1267 -77 1325 -71
rect 1459 -37 1517 -31
rect 1459 -71 1471 -37
rect 1505 -71 1517 -37
rect 1459 -77 1517 -71
rect 1651 -37 1709 -31
rect 1651 -71 1663 -37
rect 1697 -71 1709 -37
rect 1651 -77 1709 -71
rect 1843 -37 1901 -31
rect 1843 -71 1855 -37
rect 1889 -71 1901 -37
rect 1843 -77 1901 -71
rect 2035 -37 2093 -31
rect 2035 -71 2047 -37
rect 2081 -71 2093 -37
rect 2035 -77 2093 -71
rect 2227 -37 2285 -31
rect 2227 -71 2239 -37
rect 2273 -71 2285 -37
rect 2227 -77 2285 -71
rect -2423 -121 -2377 -109
rect -2423 -497 -2417 -121
rect -2383 -497 -2377 -121
rect -2423 -509 -2377 -497
rect -2327 -121 -2281 -109
rect -2327 -497 -2321 -121
rect -2287 -497 -2281 -121
rect -2327 -509 -2281 -497
rect -2231 -121 -2185 -109
rect -2231 -497 -2225 -121
rect -2191 -497 -2185 -121
rect -2231 -509 -2185 -497
rect -2135 -121 -2089 -109
rect -2135 -497 -2129 -121
rect -2095 -497 -2089 -121
rect -2135 -509 -2089 -497
rect -2039 -121 -1993 -109
rect -2039 -497 -2033 -121
rect -1999 -497 -1993 -121
rect -2039 -509 -1993 -497
rect -1943 -121 -1897 -109
rect -1943 -497 -1937 -121
rect -1903 -497 -1897 -121
rect -1943 -509 -1897 -497
rect -1847 -121 -1801 -109
rect -1847 -497 -1841 -121
rect -1807 -497 -1801 -121
rect -1847 -509 -1801 -497
rect -1751 -121 -1705 -109
rect -1751 -497 -1745 -121
rect -1711 -497 -1705 -121
rect -1751 -509 -1705 -497
rect -1655 -121 -1609 -109
rect -1655 -497 -1649 -121
rect -1615 -497 -1609 -121
rect -1655 -509 -1609 -497
rect -1559 -121 -1513 -109
rect -1559 -497 -1553 -121
rect -1519 -497 -1513 -121
rect -1559 -509 -1513 -497
rect -1463 -121 -1417 -109
rect -1463 -497 -1457 -121
rect -1423 -497 -1417 -121
rect -1463 -509 -1417 -497
rect -1367 -121 -1321 -109
rect -1367 -497 -1361 -121
rect -1327 -497 -1321 -121
rect -1367 -509 -1321 -497
rect -1271 -121 -1225 -109
rect -1271 -497 -1265 -121
rect -1231 -497 -1225 -121
rect -1271 -509 -1225 -497
rect -1175 -121 -1129 -109
rect -1175 -497 -1169 -121
rect -1135 -497 -1129 -121
rect -1175 -509 -1129 -497
rect -1079 -121 -1033 -109
rect -1079 -497 -1073 -121
rect -1039 -497 -1033 -121
rect -1079 -509 -1033 -497
rect -983 -121 -937 -109
rect -983 -497 -977 -121
rect -943 -497 -937 -121
rect -983 -509 -937 -497
rect -887 -121 -841 -109
rect -887 -497 -881 -121
rect -847 -497 -841 -121
rect -887 -509 -841 -497
rect -791 -121 -745 -109
rect -791 -497 -785 -121
rect -751 -497 -745 -121
rect -791 -509 -745 -497
rect -695 -121 -649 -109
rect -695 -497 -689 -121
rect -655 -497 -649 -121
rect -695 -509 -649 -497
rect -599 -121 -553 -109
rect -599 -497 -593 -121
rect -559 -497 -553 -121
rect -599 -509 -553 -497
rect -503 -121 -457 -109
rect -503 -497 -497 -121
rect -463 -497 -457 -121
rect -503 -509 -457 -497
rect -407 -121 -361 -109
rect -407 -497 -401 -121
rect -367 -497 -361 -121
rect -407 -509 -361 -497
rect -311 -121 -265 -109
rect -311 -497 -305 -121
rect -271 -497 -265 -121
rect -311 -509 -265 -497
rect -215 -121 -169 -109
rect -215 -497 -209 -121
rect -175 -497 -169 -121
rect -215 -509 -169 -497
rect -119 -121 -73 -109
rect -119 -497 -113 -121
rect -79 -497 -73 -121
rect -119 -509 -73 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 73 -121 119 -109
rect 73 -497 79 -121
rect 113 -497 119 -121
rect 73 -509 119 -497
rect 169 -121 215 -109
rect 169 -497 175 -121
rect 209 -497 215 -121
rect 169 -509 215 -497
rect 265 -121 311 -109
rect 265 -497 271 -121
rect 305 -497 311 -121
rect 265 -509 311 -497
rect 361 -121 407 -109
rect 361 -497 367 -121
rect 401 -497 407 -121
rect 361 -509 407 -497
rect 457 -121 503 -109
rect 457 -497 463 -121
rect 497 -497 503 -121
rect 457 -509 503 -497
rect 553 -121 599 -109
rect 553 -497 559 -121
rect 593 -497 599 -121
rect 553 -509 599 -497
rect 649 -121 695 -109
rect 649 -497 655 -121
rect 689 -497 695 -121
rect 649 -509 695 -497
rect 745 -121 791 -109
rect 745 -497 751 -121
rect 785 -497 791 -121
rect 745 -509 791 -497
rect 841 -121 887 -109
rect 841 -497 847 -121
rect 881 -497 887 -121
rect 841 -509 887 -497
rect 937 -121 983 -109
rect 937 -497 943 -121
rect 977 -497 983 -121
rect 937 -509 983 -497
rect 1033 -121 1079 -109
rect 1033 -497 1039 -121
rect 1073 -497 1079 -121
rect 1033 -509 1079 -497
rect 1129 -121 1175 -109
rect 1129 -497 1135 -121
rect 1169 -497 1175 -121
rect 1129 -509 1175 -497
rect 1225 -121 1271 -109
rect 1225 -497 1231 -121
rect 1265 -497 1271 -121
rect 1225 -509 1271 -497
rect 1321 -121 1367 -109
rect 1321 -497 1327 -121
rect 1361 -497 1367 -121
rect 1321 -509 1367 -497
rect 1417 -121 1463 -109
rect 1417 -497 1423 -121
rect 1457 -497 1463 -121
rect 1417 -509 1463 -497
rect 1513 -121 1559 -109
rect 1513 -497 1519 -121
rect 1553 -497 1559 -121
rect 1513 -509 1559 -497
rect 1609 -121 1655 -109
rect 1609 -497 1615 -121
rect 1649 -497 1655 -121
rect 1609 -509 1655 -497
rect 1705 -121 1751 -109
rect 1705 -497 1711 -121
rect 1745 -497 1751 -121
rect 1705 -509 1751 -497
rect 1801 -121 1847 -109
rect 1801 -497 1807 -121
rect 1841 -497 1847 -121
rect 1801 -509 1847 -497
rect 1897 -121 1943 -109
rect 1897 -497 1903 -121
rect 1937 -497 1943 -121
rect 1897 -509 1943 -497
rect 1993 -121 2039 -109
rect 1993 -497 1999 -121
rect 2033 -497 2039 -121
rect 1993 -509 2039 -497
rect 2089 -121 2135 -109
rect 2089 -497 2095 -121
rect 2129 -497 2135 -121
rect 2089 -509 2135 -497
rect 2185 -121 2231 -109
rect 2185 -497 2191 -121
rect 2225 -497 2231 -121
rect 2185 -509 2231 -497
rect 2281 -121 2327 -109
rect 2281 -497 2287 -121
rect 2321 -497 2327 -121
rect 2281 -509 2327 -497
rect 2377 -121 2423 -109
rect 2377 -497 2383 -121
rect 2417 -497 2423 -121
rect 2377 -509 2423 -497
rect -2285 -547 -2227 -541
rect -2285 -581 -2273 -547
rect -2239 -581 -2227 -547
rect -2285 -587 -2227 -581
rect -2093 -547 -2035 -541
rect -2093 -581 -2081 -547
rect -2047 -581 -2035 -547
rect -2093 -587 -2035 -581
rect -1901 -547 -1843 -541
rect -1901 -581 -1889 -547
rect -1855 -581 -1843 -547
rect -1901 -587 -1843 -581
rect -1709 -547 -1651 -541
rect -1709 -581 -1697 -547
rect -1663 -581 -1651 -547
rect -1709 -587 -1651 -581
rect -1517 -547 -1459 -541
rect -1517 -581 -1505 -547
rect -1471 -581 -1459 -547
rect -1517 -587 -1459 -581
rect -1325 -547 -1267 -541
rect -1325 -581 -1313 -547
rect -1279 -581 -1267 -547
rect -1325 -587 -1267 -581
rect -1133 -547 -1075 -541
rect -1133 -581 -1121 -547
rect -1087 -581 -1075 -547
rect -1133 -587 -1075 -581
rect -941 -547 -883 -541
rect -941 -581 -929 -547
rect -895 -581 -883 -547
rect -941 -587 -883 -581
rect -749 -547 -691 -541
rect -749 -581 -737 -547
rect -703 -581 -691 -547
rect -749 -587 -691 -581
rect -557 -547 -499 -541
rect -557 -581 -545 -547
rect -511 -581 -499 -547
rect -557 -587 -499 -581
rect -365 -547 -307 -541
rect -365 -581 -353 -547
rect -319 -581 -307 -547
rect -365 -587 -307 -581
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
rect 211 -547 269 -541
rect 211 -581 223 -547
rect 257 -581 269 -547
rect 211 -587 269 -581
rect 403 -547 461 -541
rect 403 -581 415 -547
rect 449 -581 461 -547
rect 403 -587 461 -581
rect 595 -547 653 -541
rect 595 -581 607 -547
rect 641 -581 653 -547
rect 595 -587 653 -581
rect 787 -547 845 -541
rect 787 -581 799 -547
rect 833 -581 845 -547
rect 787 -587 845 -581
rect 979 -547 1037 -541
rect 979 -581 991 -547
rect 1025 -581 1037 -547
rect 979 -587 1037 -581
rect 1171 -547 1229 -541
rect 1171 -581 1183 -547
rect 1217 -581 1229 -547
rect 1171 -587 1229 -581
rect 1363 -547 1421 -541
rect 1363 -581 1375 -547
rect 1409 -581 1421 -547
rect 1363 -587 1421 -581
rect 1555 -547 1613 -541
rect 1555 -581 1567 -547
rect 1601 -581 1613 -547
rect 1555 -587 1613 -581
rect 1747 -547 1805 -541
rect 1747 -581 1759 -547
rect 1793 -581 1805 -547
rect 1747 -587 1805 -581
rect 1939 -547 1997 -541
rect 1939 -581 1951 -547
rect 1985 -581 1997 -547
rect 1939 -587 1997 -581
rect 2131 -547 2189 -541
rect 2131 -581 2143 -547
rect 2177 -581 2189 -547
rect 2131 -587 2189 -581
rect 2323 -547 2381 -541
rect 2323 -581 2335 -547
rect 2369 -581 2381 -547
rect 2323 -587 2381 -581
rect -2285 -655 -2227 -649
rect -2285 -689 -2273 -655
rect -2239 -689 -2227 -655
rect -2285 -695 -2227 -689
rect -2093 -655 -2035 -649
rect -2093 -689 -2081 -655
rect -2047 -689 -2035 -655
rect -2093 -695 -2035 -689
rect -1901 -655 -1843 -649
rect -1901 -689 -1889 -655
rect -1855 -689 -1843 -655
rect -1901 -695 -1843 -689
rect -1709 -655 -1651 -649
rect -1709 -689 -1697 -655
rect -1663 -689 -1651 -655
rect -1709 -695 -1651 -689
rect -1517 -655 -1459 -649
rect -1517 -689 -1505 -655
rect -1471 -689 -1459 -655
rect -1517 -695 -1459 -689
rect -1325 -655 -1267 -649
rect -1325 -689 -1313 -655
rect -1279 -689 -1267 -655
rect -1325 -695 -1267 -689
rect -1133 -655 -1075 -649
rect -1133 -689 -1121 -655
rect -1087 -689 -1075 -655
rect -1133 -695 -1075 -689
rect -941 -655 -883 -649
rect -941 -689 -929 -655
rect -895 -689 -883 -655
rect -941 -695 -883 -689
rect -749 -655 -691 -649
rect -749 -689 -737 -655
rect -703 -689 -691 -655
rect -749 -695 -691 -689
rect -557 -655 -499 -649
rect -557 -689 -545 -655
rect -511 -689 -499 -655
rect -557 -695 -499 -689
rect -365 -655 -307 -649
rect -365 -689 -353 -655
rect -319 -689 -307 -655
rect -365 -695 -307 -689
rect -173 -655 -115 -649
rect -173 -689 -161 -655
rect -127 -689 -115 -655
rect -173 -695 -115 -689
rect 19 -655 77 -649
rect 19 -689 31 -655
rect 65 -689 77 -655
rect 19 -695 77 -689
rect 211 -655 269 -649
rect 211 -689 223 -655
rect 257 -689 269 -655
rect 211 -695 269 -689
rect 403 -655 461 -649
rect 403 -689 415 -655
rect 449 -689 461 -655
rect 403 -695 461 -689
rect 595 -655 653 -649
rect 595 -689 607 -655
rect 641 -689 653 -655
rect 595 -695 653 -689
rect 787 -655 845 -649
rect 787 -689 799 -655
rect 833 -689 845 -655
rect 787 -695 845 -689
rect 979 -655 1037 -649
rect 979 -689 991 -655
rect 1025 -689 1037 -655
rect 979 -695 1037 -689
rect 1171 -655 1229 -649
rect 1171 -689 1183 -655
rect 1217 -689 1229 -655
rect 1171 -695 1229 -689
rect 1363 -655 1421 -649
rect 1363 -689 1375 -655
rect 1409 -689 1421 -655
rect 1363 -695 1421 -689
rect 1555 -655 1613 -649
rect 1555 -689 1567 -655
rect 1601 -689 1613 -655
rect 1555 -695 1613 -689
rect 1747 -655 1805 -649
rect 1747 -689 1759 -655
rect 1793 -689 1805 -655
rect 1747 -695 1805 -689
rect 1939 -655 1997 -649
rect 1939 -689 1951 -655
rect 1985 -689 1997 -655
rect 1939 -695 1997 -689
rect 2131 -655 2189 -649
rect 2131 -689 2143 -655
rect 2177 -689 2189 -655
rect 2131 -695 2189 -689
rect 2323 -655 2381 -649
rect 2323 -689 2335 -655
rect 2369 -689 2381 -655
rect 2323 -695 2381 -689
rect -2423 -739 -2377 -727
rect -2423 -1115 -2417 -739
rect -2383 -1115 -2377 -739
rect -2423 -1127 -2377 -1115
rect -2327 -739 -2281 -727
rect -2327 -1115 -2321 -739
rect -2287 -1115 -2281 -739
rect -2327 -1127 -2281 -1115
rect -2231 -739 -2185 -727
rect -2231 -1115 -2225 -739
rect -2191 -1115 -2185 -739
rect -2231 -1127 -2185 -1115
rect -2135 -739 -2089 -727
rect -2135 -1115 -2129 -739
rect -2095 -1115 -2089 -739
rect -2135 -1127 -2089 -1115
rect -2039 -739 -1993 -727
rect -2039 -1115 -2033 -739
rect -1999 -1115 -1993 -739
rect -2039 -1127 -1993 -1115
rect -1943 -739 -1897 -727
rect -1943 -1115 -1937 -739
rect -1903 -1115 -1897 -739
rect -1943 -1127 -1897 -1115
rect -1847 -739 -1801 -727
rect -1847 -1115 -1841 -739
rect -1807 -1115 -1801 -739
rect -1847 -1127 -1801 -1115
rect -1751 -739 -1705 -727
rect -1751 -1115 -1745 -739
rect -1711 -1115 -1705 -739
rect -1751 -1127 -1705 -1115
rect -1655 -739 -1609 -727
rect -1655 -1115 -1649 -739
rect -1615 -1115 -1609 -739
rect -1655 -1127 -1609 -1115
rect -1559 -739 -1513 -727
rect -1559 -1115 -1553 -739
rect -1519 -1115 -1513 -739
rect -1559 -1127 -1513 -1115
rect -1463 -739 -1417 -727
rect -1463 -1115 -1457 -739
rect -1423 -1115 -1417 -739
rect -1463 -1127 -1417 -1115
rect -1367 -739 -1321 -727
rect -1367 -1115 -1361 -739
rect -1327 -1115 -1321 -739
rect -1367 -1127 -1321 -1115
rect -1271 -739 -1225 -727
rect -1271 -1115 -1265 -739
rect -1231 -1115 -1225 -739
rect -1271 -1127 -1225 -1115
rect -1175 -739 -1129 -727
rect -1175 -1115 -1169 -739
rect -1135 -1115 -1129 -739
rect -1175 -1127 -1129 -1115
rect -1079 -739 -1033 -727
rect -1079 -1115 -1073 -739
rect -1039 -1115 -1033 -739
rect -1079 -1127 -1033 -1115
rect -983 -739 -937 -727
rect -983 -1115 -977 -739
rect -943 -1115 -937 -739
rect -983 -1127 -937 -1115
rect -887 -739 -841 -727
rect -887 -1115 -881 -739
rect -847 -1115 -841 -739
rect -887 -1127 -841 -1115
rect -791 -739 -745 -727
rect -791 -1115 -785 -739
rect -751 -1115 -745 -739
rect -791 -1127 -745 -1115
rect -695 -739 -649 -727
rect -695 -1115 -689 -739
rect -655 -1115 -649 -739
rect -695 -1127 -649 -1115
rect -599 -739 -553 -727
rect -599 -1115 -593 -739
rect -559 -1115 -553 -739
rect -599 -1127 -553 -1115
rect -503 -739 -457 -727
rect -503 -1115 -497 -739
rect -463 -1115 -457 -739
rect -503 -1127 -457 -1115
rect -407 -739 -361 -727
rect -407 -1115 -401 -739
rect -367 -1115 -361 -739
rect -407 -1127 -361 -1115
rect -311 -739 -265 -727
rect -311 -1115 -305 -739
rect -271 -1115 -265 -739
rect -311 -1127 -265 -1115
rect -215 -739 -169 -727
rect -215 -1115 -209 -739
rect -175 -1115 -169 -739
rect -215 -1127 -169 -1115
rect -119 -739 -73 -727
rect -119 -1115 -113 -739
rect -79 -1115 -73 -739
rect -119 -1127 -73 -1115
rect -23 -739 23 -727
rect -23 -1115 -17 -739
rect 17 -1115 23 -739
rect -23 -1127 23 -1115
rect 73 -739 119 -727
rect 73 -1115 79 -739
rect 113 -1115 119 -739
rect 73 -1127 119 -1115
rect 169 -739 215 -727
rect 169 -1115 175 -739
rect 209 -1115 215 -739
rect 169 -1127 215 -1115
rect 265 -739 311 -727
rect 265 -1115 271 -739
rect 305 -1115 311 -739
rect 265 -1127 311 -1115
rect 361 -739 407 -727
rect 361 -1115 367 -739
rect 401 -1115 407 -739
rect 361 -1127 407 -1115
rect 457 -739 503 -727
rect 457 -1115 463 -739
rect 497 -1115 503 -739
rect 457 -1127 503 -1115
rect 553 -739 599 -727
rect 553 -1115 559 -739
rect 593 -1115 599 -739
rect 553 -1127 599 -1115
rect 649 -739 695 -727
rect 649 -1115 655 -739
rect 689 -1115 695 -739
rect 649 -1127 695 -1115
rect 745 -739 791 -727
rect 745 -1115 751 -739
rect 785 -1115 791 -739
rect 745 -1127 791 -1115
rect 841 -739 887 -727
rect 841 -1115 847 -739
rect 881 -1115 887 -739
rect 841 -1127 887 -1115
rect 937 -739 983 -727
rect 937 -1115 943 -739
rect 977 -1115 983 -739
rect 937 -1127 983 -1115
rect 1033 -739 1079 -727
rect 1033 -1115 1039 -739
rect 1073 -1115 1079 -739
rect 1033 -1127 1079 -1115
rect 1129 -739 1175 -727
rect 1129 -1115 1135 -739
rect 1169 -1115 1175 -739
rect 1129 -1127 1175 -1115
rect 1225 -739 1271 -727
rect 1225 -1115 1231 -739
rect 1265 -1115 1271 -739
rect 1225 -1127 1271 -1115
rect 1321 -739 1367 -727
rect 1321 -1115 1327 -739
rect 1361 -1115 1367 -739
rect 1321 -1127 1367 -1115
rect 1417 -739 1463 -727
rect 1417 -1115 1423 -739
rect 1457 -1115 1463 -739
rect 1417 -1127 1463 -1115
rect 1513 -739 1559 -727
rect 1513 -1115 1519 -739
rect 1553 -1115 1559 -739
rect 1513 -1127 1559 -1115
rect 1609 -739 1655 -727
rect 1609 -1115 1615 -739
rect 1649 -1115 1655 -739
rect 1609 -1127 1655 -1115
rect 1705 -739 1751 -727
rect 1705 -1115 1711 -739
rect 1745 -1115 1751 -739
rect 1705 -1127 1751 -1115
rect 1801 -739 1847 -727
rect 1801 -1115 1807 -739
rect 1841 -1115 1847 -739
rect 1801 -1127 1847 -1115
rect 1897 -739 1943 -727
rect 1897 -1115 1903 -739
rect 1937 -1115 1943 -739
rect 1897 -1127 1943 -1115
rect 1993 -739 2039 -727
rect 1993 -1115 1999 -739
rect 2033 -1115 2039 -739
rect 1993 -1127 2039 -1115
rect 2089 -739 2135 -727
rect 2089 -1115 2095 -739
rect 2129 -1115 2135 -739
rect 2089 -1127 2135 -1115
rect 2185 -739 2231 -727
rect 2185 -1115 2191 -739
rect 2225 -1115 2231 -739
rect 2185 -1127 2231 -1115
rect 2281 -739 2327 -727
rect 2281 -1115 2287 -739
rect 2321 -1115 2327 -739
rect 2281 -1127 2327 -1115
rect 2377 -739 2423 -727
rect 2377 -1115 2383 -739
rect 2417 -1115 2423 -739
rect 2377 -1127 2423 -1115
rect -2381 -1165 -2323 -1159
rect -2381 -1199 -2369 -1165
rect -2335 -1199 -2323 -1165
rect -2381 -1205 -2323 -1199
rect -2189 -1165 -2131 -1159
rect -2189 -1199 -2177 -1165
rect -2143 -1199 -2131 -1165
rect -2189 -1205 -2131 -1199
rect -1997 -1165 -1939 -1159
rect -1997 -1199 -1985 -1165
rect -1951 -1199 -1939 -1165
rect -1997 -1205 -1939 -1199
rect -1805 -1165 -1747 -1159
rect -1805 -1199 -1793 -1165
rect -1759 -1199 -1747 -1165
rect -1805 -1205 -1747 -1199
rect -1613 -1165 -1555 -1159
rect -1613 -1199 -1601 -1165
rect -1567 -1199 -1555 -1165
rect -1613 -1205 -1555 -1199
rect -1421 -1165 -1363 -1159
rect -1421 -1199 -1409 -1165
rect -1375 -1199 -1363 -1165
rect -1421 -1205 -1363 -1199
rect -1229 -1165 -1171 -1159
rect -1229 -1199 -1217 -1165
rect -1183 -1199 -1171 -1165
rect -1229 -1205 -1171 -1199
rect -1037 -1165 -979 -1159
rect -1037 -1199 -1025 -1165
rect -991 -1199 -979 -1165
rect -1037 -1205 -979 -1199
rect -845 -1165 -787 -1159
rect -845 -1199 -833 -1165
rect -799 -1199 -787 -1165
rect -845 -1205 -787 -1199
rect -653 -1165 -595 -1159
rect -653 -1199 -641 -1165
rect -607 -1199 -595 -1165
rect -653 -1205 -595 -1199
rect -461 -1165 -403 -1159
rect -461 -1199 -449 -1165
rect -415 -1199 -403 -1165
rect -461 -1205 -403 -1199
rect -269 -1165 -211 -1159
rect -269 -1199 -257 -1165
rect -223 -1199 -211 -1165
rect -269 -1205 -211 -1199
rect -77 -1165 -19 -1159
rect -77 -1199 -65 -1165
rect -31 -1199 -19 -1165
rect -77 -1205 -19 -1199
rect 115 -1165 173 -1159
rect 115 -1199 127 -1165
rect 161 -1199 173 -1165
rect 115 -1205 173 -1199
rect 307 -1165 365 -1159
rect 307 -1199 319 -1165
rect 353 -1199 365 -1165
rect 307 -1205 365 -1199
rect 499 -1165 557 -1159
rect 499 -1199 511 -1165
rect 545 -1199 557 -1165
rect 499 -1205 557 -1199
rect 691 -1165 749 -1159
rect 691 -1199 703 -1165
rect 737 -1199 749 -1165
rect 691 -1205 749 -1199
rect 883 -1165 941 -1159
rect 883 -1199 895 -1165
rect 929 -1199 941 -1165
rect 883 -1205 941 -1199
rect 1075 -1165 1133 -1159
rect 1075 -1199 1087 -1165
rect 1121 -1199 1133 -1165
rect 1075 -1205 1133 -1199
rect 1267 -1165 1325 -1159
rect 1267 -1199 1279 -1165
rect 1313 -1199 1325 -1165
rect 1267 -1205 1325 -1199
rect 1459 -1165 1517 -1159
rect 1459 -1199 1471 -1165
rect 1505 -1199 1517 -1165
rect 1459 -1205 1517 -1199
rect 1651 -1165 1709 -1159
rect 1651 -1199 1663 -1165
rect 1697 -1199 1709 -1165
rect 1651 -1205 1709 -1199
rect 1843 -1165 1901 -1159
rect 1843 -1199 1855 -1165
rect 1889 -1199 1901 -1165
rect 1843 -1205 1901 -1199
rect 2035 -1165 2093 -1159
rect 2035 -1199 2047 -1165
rect 2081 -1199 2093 -1165
rect 2035 -1205 2093 -1199
rect 2227 -1165 2285 -1159
rect 2227 -1199 2239 -1165
rect 2273 -1199 2285 -1165
rect 2227 -1205 2285 -1199
<< properties >>
string FIXED_BBOX -2514 -1284 2514 1284
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 4 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
