magic
tech sky130A
magscale 1 2
timestamp 1646400034
<< error_p >>
rect -78 181 -20 187
rect 118 181 176 187
rect -78 147 -66 181
rect 118 147 130 181
rect -78 141 -20 147
rect 118 141 176 147
rect -176 -147 -118 -141
rect 20 -147 78 -141
rect -176 -181 -164 -147
rect 20 -181 32 -147
rect -176 -187 -118 -181
rect 20 -187 78 -181
<< nwell >>
rect -363 -319 363 319
<< pmos >>
rect -167 -100 -127 100
rect -69 -100 -29 100
rect 29 -100 69 100
rect 127 -100 167 100
<< pdiff >>
rect -225 88 -167 100
rect -225 -88 -213 88
rect -179 -88 -167 88
rect -225 -100 -167 -88
rect -127 88 -69 100
rect -127 -88 -115 88
rect -81 -88 -69 88
rect -127 -100 -69 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 69 88 127 100
rect 69 -88 81 88
rect 115 -88 127 88
rect 69 -100 127 -88
rect 167 88 225 100
rect 167 -88 179 88
rect 213 -88 225 88
rect 167 -100 225 -88
<< pdiffc >>
rect -213 -88 -179 88
rect -115 -88 -81 88
rect -17 -88 17 88
rect 81 -88 115 88
rect 179 -88 213 88
<< nsubdiff >>
rect -327 249 -231 283
rect 231 249 327 283
rect -327 187 -293 249
rect 293 187 327 249
rect -327 -249 -293 -187
rect 293 -249 327 -187
rect -327 -283 -231 -249
rect 231 -283 327 -249
<< nsubdiffcont >>
rect -231 249 231 283
rect -327 -187 -293 187
rect 293 -187 327 187
rect -231 -283 231 -249
<< poly >>
rect -82 181 -16 197
rect -82 147 -66 181
rect -32 147 -16 181
rect -82 131 -16 147
rect 114 181 180 197
rect 114 147 130 181
rect 164 147 180 181
rect 114 131 180 147
rect -167 100 -127 126
rect -69 100 -29 131
rect 29 100 69 126
rect 127 100 167 131
rect -167 -131 -127 -100
rect -69 -126 -29 -100
rect 29 -131 69 -100
rect 127 -126 167 -100
rect -180 -147 -114 -131
rect -180 -181 -164 -147
rect -130 -181 -114 -147
rect -180 -197 -114 -181
rect 16 -147 82 -131
rect 16 -181 32 -147
rect 66 -181 82 -147
rect 16 -197 82 -181
<< polycont >>
rect -66 147 -32 181
rect 130 147 164 181
rect -164 -181 -130 -147
rect 32 -181 66 -147
<< locali >>
rect -327 249 -231 283
rect 231 249 327 283
rect -327 187 -293 249
rect 293 187 327 249
rect -82 147 -66 181
rect -32 147 -16 181
rect 114 147 130 181
rect 164 147 180 181
rect -213 88 -179 104
rect -213 -104 -179 -88
rect -115 88 -81 104
rect -115 -104 -81 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 81 88 115 104
rect 81 -104 115 -88
rect 179 88 213 104
rect 179 -104 213 -88
rect -180 -181 -164 -147
rect -130 -181 -114 -147
rect 16 -181 32 -147
rect 66 -181 82 -147
rect -327 -249 -293 -187
rect 293 -249 327 -187
rect -327 -283 -231 -249
rect 231 -283 327 -249
<< viali >>
rect -66 147 -32 181
rect 130 147 164 181
rect -213 -88 -179 88
rect -115 -88 -81 88
rect -17 -88 17 88
rect 81 -88 115 88
rect 179 -88 213 88
rect -164 -181 -130 -147
rect 32 -181 66 -147
<< metal1 >>
rect -78 181 -20 187
rect -78 147 -66 181
rect -32 147 -20 181
rect -78 141 -20 147
rect 118 181 176 187
rect 118 147 130 181
rect 164 147 176 181
rect 118 141 176 147
rect -219 88 -173 100
rect -219 -88 -213 88
rect -179 -88 -173 88
rect -219 -100 -173 -88
rect -121 88 -75 100
rect -121 -88 -115 88
rect -81 -88 -75 88
rect -121 -100 -75 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 75 88 121 100
rect 75 -88 81 88
rect 115 -88 121 88
rect 75 -100 121 -88
rect 173 88 219 100
rect 173 -88 179 88
rect 213 -88 219 88
rect 173 -100 219 -88
rect -176 -147 -118 -141
rect -176 -181 -164 -147
rect -130 -181 -118 -147
rect -176 -187 -118 -181
rect 20 -147 78 -141
rect 20 -181 32 -147
rect 66 -181 78 -147
rect 20 -187 78 -181
<< properties >>
string FIXED_BBOX -310 -266 310 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.2 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
