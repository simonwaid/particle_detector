magic
tech sky130A
magscale 1 2
timestamp 1645462850
<< pwell >>
rect -3312 -2137 3312 2137
<< nmos >>
rect -3116 1127 -1916 1927
rect -1858 1127 -658 1927
rect -600 1127 600 1927
rect 658 1127 1858 1927
rect 1916 1127 3116 1927
rect -3116 109 -1916 909
rect -1858 109 -658 909
rect -600 109 600 909
rect 658 109 1858 909
rect 1916 109 3116 909
rect -3116 -909 -1916 -109
rect -1858 -909 -658 -109
rect -600 -909 600 -109
rect 658 -909 1858 -109
rect 1916 -909 3116 -109
rect -3116 -1927 -1916 -1127
rect -1858 -1927 -658 -1127
rect -600 -1927 600 -1127
rect 658 -1927 1858 -1127
rect 1916 -1927 3116 -1127
<< ndiff >>
rect -3174 1915 -3116 1927
rect -3174 1139 -3162 1915
rect -3128 1139 -3116 1915
rect -3174 1127 -3116 1139
rect -1916 1915 -1858 1927
rect -1916 1139 -1904 1915
rect -1870 1139 -1858 1915
rect -1916 1127 -1858 1139
rect -658 1915 -600 1927
rect -658 1139 -646 1915
rect -612 1139 -600 1915
rect -658 1127 -600 1139
rect 600 1915 658 1927
rect 600 1139 612 1915
rect 646 1139 658 1915
rect 600 1127 658 1139
rect 1858 1915 1916 1927
rect 1858 1139 1870 1915
rect 1904 1139 1916 1915
rect 1858 1127 1916 1139
rect 3116 1915 3174 1927
rect 3116 1139 3128 1915
rect 3162 1139 3174 1915
rect 3116 1127 3174 1139
rect -3174 897 -3116 909
rect -3174 121 -3162 897
rect -3128 121 -3116 897
rect -3174 109 -3116 121
rect -1916 897 -1858 909
rect -1916 121 -1904 897
rect -1870 121 -1858 897
rect -1916 109 -1858 121
rect -658 897 -600 909
rect -658 121 -646 897
rect -612 121 -600 897
rect -658 109 -600 121
rect 600 897 658 909
rect 600 121 612 897
rect 646 121 658 897
rect 600 109 658 121
rect 1858 897 1916 909
rect 1858 121 1870 897
rect 1904 121 1916 897
rect 1858 109 1916 121
rect 3116 897 3174 909
rect 3116 121 3128 897
rect 3162 121 3174 897
rect 3116 109 3174 121
rect -3174 -121 -3116 -109
rect -3174 -897 -3162 -121
rect -3128 -897 -3116 -121
rect -3174 -909 -3116 -897
rect -1916 -121 -1858 -109
rect -1916 -897 -1904 -121
rect -1870 -897 -1858 -121
rect -1916 -909 -1858 -897
rect -658 -121 -600 -109
rect -658 -897 -646 -121
rect -612 -897 -600 -121
rect -658 -909 -600 -897
rect 600 -121 658 -109
rect 600 -897 612 -121
rect 646 -897 658 -121
rect 600 -909 658 -897
rect 1858 -121 1916 -109
rect 1858 -897 1870 -121
rect 1904 -897 1916 -121
rect 1858 -909 1916 -897
rect 3116 -121 3174 -109
rect 3116 -897 3128 -121
rect 3162 -897 3174 -121
rect 3116 -909 3174 -897
rect -3174 -1139 -3116 -1127
rect -3174 -1915 -3162 -1139
rect -3128 -1915 -3116 -1139
rect -3174 -1927 -3116 -1915
rect -1916 -1139 -1858 -1127
rect -1916 -1915 -1904 -1139
rect -1870 -1915 -1858 -1139
rect -1916 -1927 -1858 -1915
rect -658 -1139 -600 -1127
rect -658 -1915 -646 -1139
rect -612 -1915 -600 -1139
rect -658 -1927 -600 -1915
rect 600 -1139 658 -1127
rect 600 -1915 612 -1139
rect 646 -1915 658 -1139
rect 600 -1927 658 -1915
rect 1858 -1139 1916 -1127
rect 1858 -1915 1870 -1139
rect 1904 -1915 1916 -1139
rect 1858 -1927 1916 -1915
rect 3116 -1139 3174 -1127
rect 3116 -1915 3128 -1139
rect 3162 -1915 3174 -1139
rect 3116 -1927 3174 -1915
<< ndiffc >>
rect -3162 1139 -3128 1915
rect -1904 1139 -1870 1915
rect -646 1139 -612 1915
rect 612 1139 646 1915
rect 1870 1139 1904 1915
rect 3128 1139 3162 1915
rect -3162 121 -3128 897
rect -1904 121 -1870 897
rect -646 121 -612 897
rect 612 121 646 897
rect 1870 121 1904 897
rect 3128 121 3162 897
rect -3162 -897 -3128 -121
rect -1904 -897 -1870 -121
rect -646 -897 -612 -121
rect 612 -897 646 -121
rect 1870 -897 1904 -121
rect 3128 -897 3162 -121
rect -3162 -1915 -3128 -1139
rect -1904 -1915 -1870 -1139
rect -646 -1915 -612 -1139
rect 612 -1915 646 -1139
rect 1870 -1915 1904 -1139
rect 3128 -1915 3162 -1139
<< psubdiff >>
rect -3276 2067 -3180 2101
rect 3180 2067 3276 2101
rect -3276 2005 -3242 2067
rect 3242 2005 3276 2067
rect -3276 -2067 -3242 -2005
rect 3242 -2067 3276 -2005
rect -3276 -2101 -3180 -2067
rect 3180 -2101 3276 -2067
<< psubdiffcont >>
rect -3180 2067 3180 2101
rect -3276 -2005 -3242 2005
rect 3242 -2005 3276 2005
rect -3180 -2101 3180 -2067
<< poly >>
rect -3116 1999 -1916 2015
rect -3116 1965 -3100 1999
rect -1932 1965 -1916 1999
rect -3116 1927 -1916 1965
rect -1858 1999 -658 2015
rect -1858 1965 -1842 1999
rect -674 1965 -658 1999
rect -1858 1927 -658 1965
rect -600 1999 600 2015
rect -600 1965 -584 1999
rect 584 1965 600 1999
rect -600 1927 600 1965
rect 658 1999 1858 2015
rect 658 1965 674 1999
rect 1842 1965 1858 1999
rect 658 1927 1858 1965
rect 1916 1999 3116 2015
rect 1916 1965 1932 1999
rect 3100 1965 3116 1999
rect 1916 1927 3116 1965
rect -3116 1089 -1916 1127
rect -3116 1055 -3100 1089
rect -1932 1055 -1916 1089
rect -3116 1039 -1916 1055
rect -1858 1089 -658 1127
rect -1858 1055 -1842 1089
rect -674 1055 -658 1089
rect -1858 1039 -658 1055
rect -600 1089 600 1127
rect -600 1055 -584 1089
rect 584 1055 600 1089
rect -600 1039 600 1055
rect 658 1089 1858 1127
rect 658 1055 674 1089
rect 1842 1055 1858 1089
rect 658 1039 1858 1055
rect 1916 1089 3116 1127
rect 1916 1055 1932 1089
rect 3100 1055 3116 1089
rect 1916 1039 3116 1055
rect -3116 981 -1916 997
rect -3116 947 -3100 981
rect -1932 947 -1916 981
rect -3116 909 -1916 947
rect -1858 981 -658 997
rect -1858 947 -1842 981
rect -674 947 -658 981
rect -1858 909 -658 947
rect -600 981 600 997
rect -600 947 -584 981
rect 584 947 600 981
rect -600 909 600 947
rect 658 981 1858 997
rect 658 947 674 981
rect 1842 947 1858 981
rect 658 909 1858 947
rect 1916 981 3116 997
rect 1916 947 1932 981
rect 3100 947 3116 981
rect 1916 909 3116 947
rect -3116 71 -1916 109
rect -3116 37 -3100 71
rect -1932 37 -1916 71
rect -3116 21 -1916 37
rect -1858 71 -658 109
rect -1858 37 -1842 71
rect -674 37 -658 71
rect -1858 21 -658 37
rect -600 71 600 109
rect -600 37 -584 71
rect 584 37 600 71
rect -600 21 600 37
rect 658 71 1858 109
rect 658 37 674 71
rect 1842 37 1858 71
rect 658 21 1858 37
rect 1916 71 3116 109
rect 1916 37 1932 71
rect 3100 37 3116 71
rect 1916 21 3116 37
rect -3116 -37 -1916 -21
rect -3116 -71 -3100 -37
rect -1932 -71 -1916 -37
rect -3116 -109 -1916 -71
rect -1858 -37 -658 -21
rect -1858 -71 -1842 -37
rect -674 -71 -658 -37
rect -1858 -109 -658 -71
rect -600 -37 600 -21
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -600 -109 600 -71
rect 658 -37 1858 -21
rect 658 -71 674 -37
rect 1842 -71 1858 -37
rect 658 -109 1858 -71
rect 1916 -37 3116 -21
rect 1916 -71 1932 -37
rect 3100 -71 3116 -37
rect 1916 -109 3116 -71
rect -3116 -947 -1916 -909
rect -3116 -981 -3100 -947
rect -1932 -981 -1916 -947
rect -3116 -997 -1916 -981
rect -1858 -947 -658 -909
rect -1858 -981 -1842 -947
rect -674 -981 -658 -947
rect -1858 -997 -658 -981
rect -600 -947 600 -909
rect -600 -981 -584 -947
rect 584 -981 600 -947
rect -600 -997 600 -981
rect 658 -947 1858 -909
rect 658 -981 674 -947
rect 1842 -981 1858 -947
rect 658 -997 1858 -981
rect 1916 -947 3116 -909
rect 1916 -981 1932 -947
rect 3100 -981 3116 -947
rect 1916 -997 3116 -981
rect -3116 -1055 -1916 -1039
rect -3116 -1089 -3100 -1055
rect -1932 -1089 -1916 -1055
rect -3116 -1127 -1916 -1089
rect -1858 -1055 -658 -1039
rect -1858 -1089 -1842 -1055
rect -674 -1089 -658 -1055
rect -1858 -1127 -658 -1089
rect -600 -1055 600 -1039
rect -600 -1089 -584 -1055
rect 584 -1089 600 -1055
rect -600 -1127 600 -1089
rect 658 -1055 1858 -1039
rect 658 -1089 674 -1055
rect 1842 -1089 1858 -1055
rect 658 -1127 1858 -1089
rect 1916 -1055 3116 -1039
rect 1916 -1089 1932 -1055
rect 3100 -1089 3116 -1055
rect 1916 -1127 3116 -1089
rect -3116 -1965 -1916 -1927
rect -3116 -1999 -3100 -1965
rect -1932 -1999 -1916 -1965
rect -3116 -2015 -1916 -1999
rect -1858 -1965 -658 -1927
rect -1858 -1999 -1842 -1965
rect -674 -1999 -658 -1965
rect -1858 -2015 -658 -1999
rect -600 -1965 600 -1927
rect -600 -1999 -584 -1965
rect 584 -1999 600 -1965
rect -600 -2015 600 -1999
rect 658 -1965 1858 -1927
rect 658 -1999 674 -1965
rect 1842 -1999 1858 -1965
rect 658 -2015 1858 -1999
rect 1916 -1965 3116 -1927
rect 1916 -1999 1932 -1965
rect 3100 -1999 3116 -1965
rect 1916 -2015 3116 -1999
<< polycont >>
rect -3100 1965 -1932 1999
rect -1842 1965 -674 1999
rect -584 1965 584 1999
rect 674 1965 1842 1999
rect 1932 1965 3100 1999
rect -3100 1055 -1932 1089
rect -1842 1055 -674 1089
rect -584 1055 584 1089
rect 674 1055 1842 1089
rect 1932 1055 3100 1089
rect -3100 947 -1932 981
rect -1842 947 -674 981
rect -584 947 584 981
rect 674 947 1842 981
rect 1932 947 3100 981
rect -3100 37 -1932 71
rect -1842 37 -674 71
rect -584 37 584 71
rect 674 37 1842 71
rect 1932 37 3100 71
rect -3100 -71 -1932 -37
rect -1842 -71 -674 -37
rect -584 -71 584 -37
rect 674 -71 1842 -37
rect 1932 -71 3100 -37
rect -3100 -981 -1932 -947
rect -1842 -981 -674 -947
rect -584 -981 584 -947
rect 674 -981 1842 -947
rect 1932 -981 3100 -947
rect -3100 -1089 -1932 -1055
rect -1842 -1089 -674 -1055
rect -584 -1089 584 -1055
rect 674 -1089 1842 -1055
rect 1932 -1089 3100 -1055
rect -3100 -1999 -1932 -1965
rect -1842 -1999 -674 -1965
rect -584 -1999 584 -1965
rect 674 -1999 1842 -1965
rect 1932 -1999 3100 -1965
<< locali >>
rect -3276 2067 -3180 2101
rect 3180 2067 3276 2101
rect -3276 2005 -3242 2067
rect 3242 2005 3276 2067
rect -3116 1965 -3100 1999
rect -1932 1965 -1916 1999
rect -1858 1965 -1842 1999
rect -674 1965 -658 1999
rect -600 1965 -584 1999
rect 584 1965 600 1999
rect 658 1965 674 1999
rect 1842 1965 1858 1999
rect 1916 1965 1932 1999
rect 3100 1965 3116 1999
rect -3162 1915 -3128 1931
rect -3162 1123 -3128 1139
rect -1904 1915 -1870 1931
rect -1904 1123 -1870 1139
rect -646 1915 -612 1931
rect -646 1123 -612 1139
rect 612 1915 646 1931
rect 612 1123 646 1139
rect 1870 1915 1904 1931
rect 1870 1123 1904 1139
rect 3128 1915 3162 1931
rect 3128 1123 3162 1139
rect -3116 1055 -3100 1089
rect -1932 1055 -1916 1089
rect -1858 1055 -1842 1089
rect -674 1055 -658 1089
rect -600 1055 -584 1089
rect 584 1055 600 1089
rect 658 1055 674 1089
rect 1842 1055 1858 1089
rect 1916 1055 1932 1089
rect 3100 1055 3116 1089
rect -3116 947 -3100 981
rect -1932 947 -1916 981
rect -1858 947 -1842 981
rect -674 947 -658 981
rect -600 947 -584 981
rect 584 947 600 981
rect 658 947 674 981
rect 1842 947 1858 981
rect 1916 947 1932 981
rect 3100 947 3116 981
rect -3162 897 -3128 913
rect -3162 105 -3128 121
rect -1904 897 -1870 913
rect -1904 105 -1870 121
rect -646 897 -612 913
rect -646 105 -612 121
rect 612 897 646 913
rect 612 105 646 121
rect 1870 897 1904 913
rect 1870 105 1904 121
rect 3128 897 3162 913
rect 3128 105 3162 121
rect -3116 37 -3100 71
rect -1932 37 -1916 71
rect -1858 37 -1842 71
rect -674 37 -658 71
rect -600 37 -584 71
rect 584 37 600 71
rect 658 37 674 71
rect 1842 37 1858 71
rect 1916 37 1932 71
rect 3100 37 3116 71
rect -3116 -71 -3100 -37
rect -1932 -71 -1916 -37
rect -1858 -71 -1842 -37
rect -674 -71 -658 -37
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect 658 -71 674 -37
rect 1842 -71 1858 -37
rect 1916 -71 1932 -37
rect 3100 -71 3116 -37
rect -3162 -121 -3128 -105
rect -3162 -913 -3128 -897
rect -1904 -121 -1870 -105
rect -1904 -913 -1870 -897
rect -646 -121 -612 -105
rect -646 -913 -612 -897
rect 612 -121 646 -105
rect 612 -913 646 -897
rect 1870 -121 1904 -105
rect 1870 -913 1904 -897
rect 3128 -121 3162 -105
rect 3128 -913 3162 -897
rect -3116 -981 -3100 -947
rect -1932 -981 -1916 -947
rect -1858 -981 -1842 -947
rect -674 -981 -658 -947
rect -600 -981 -584 -947
rect 584 -981 600 -947
rect 658 -981 674 -947
rect 1842 -981 1858 -947
rect 1916 -981 1932 -947
rect 3100 -981 3116 -947
rect -3116 -1089 -3100 -1055
rect -1932 -1089 -1916 -1055
rect -1858 -1089 -1842 -1055
rect -674 -1089 -658 -1055
rect -600 -1089 -584 -1055
rect 584 -1089 600 -1055
rect 658 -1089 674 -1055
rect 1842 -1089 1858 -1055
rect 1916 -1089 1932 -1055
rect 3100 -1089 3116 -1055
rect -3162 -1139 -3128 -1123
rect -3162 -1931 -3128 -1915
rect -1904 -1139 -1870 -1123
rect -1904 -1931 -1870 -1915
rect -646 -1139 -612 -1123
rect -646 -1931 -612 -1915
rect 612 -1139 646 -1123
rect 612 -1931 646 -1915
rect 1870 -1139 1904 -1123
rect 1870 -1931 1904 -1915
rect 3128 -1139 3162 -1123
rect 3128 -1931 3162 -1915
rect -3116 -1999 -3100 -1965
rect -1932 -1999 -1916 -1965
rect -1858 -1999 -1842 -1965
rect -674 -1999 -658 -1965
rect -600 -1999 -584 -1965
rect 584 -1999 600 -1965
rect 658 -1999 674 -1965
rect 1842 -1999 1858 -1965
rect 1916 -1999 1932 -1965
rect 3100 -1999 3116 -1965
rect -3276 -2067 -3242 -2005
rect 3242 -2067 3276 -2005
rect -3276 -2101 -3180 -2067
rect 3180 -2101 3276 -2067
<< viali >>
rect -3100 1965 -1932 1999
rect -1842 1965 -674 1999
rect -584 1965 584 1999
rect 674 1965 1842 1999
rect 1932 1965 3100 1999
rect -3162 1139 -3128 1915
rect -1904 1139 -1870 1915
rect -646 1139 -612 1915
rect 612 1139 646 1915
rect 1870 1139 1904 1915
rect 3128 1139 3162 1915
rect -3100 1055 -1932 1089
rect -1842 1055 -674 1089
rect -584 1055 584 1089
rect 674 1055 1842 1089
rect 1932 1055 3100 1089
rect -3100 947 -1932 981
rect -1842 947 -674 981
rect -584 947 584 981
rect 674 947 1842 981
rect 1932 947 3100 981
rect -3162 121 -3128 897
rect -1904 121 -1870 897
rect -646 121 -612 897
rect 612 121 646 897
rect 1870 121 1904 897
rect 3128 121 3162 897
rect -3100 37 -1932 71
rect -1842 37 -674 71
rect -584 37 584 71
rect 674 37 1842 71
rect 1932 37 3100 71
rect -3100 -71 -1932 -37
rect -1842 -71 -674 -37
rect -584 -71 584 -37
rect 674 -71 1842 -37
rect 1932 -71 3100 -37
rect -3162 -897 -3128 -121
rect -1904 -897 -1870 -121
rect -646 -897 -612 -121
rect 612 -897 646 -121
rect 1870 -897 1904 -121
rect 3128 -897 3162 -121
rect -3100 -981 -1932 -947
rect -1842 -981 -674 -947
rect -584 -981 584 -947
rect 674 -981 1842 -947
rect 1932 -981 3100 -947
rect -3100 -1089 -1932 -1055
rect -1842 -1089 -674 -1055
rect -584 -1089 584 -1055
rect 674 -1089 1842 -1055
rect 1932 -1089 3100 -1055
rect -3162 -1915 -3128 -1139
rect -1904 -1915 -1870 -1139
rect -646 -1915 -612 -1139
rect 612 -1915 646 -1139
rect 1870 -1915 1904 -1139
rect 3128 -1915 3162 -1139
rect -3100 -1999 -1932 -1965
rect -1842 -1999 -674 -1965
rect -584 -1999 584 -1965
rect 674 -1999 1842 -1965
rect 1932 -1999 3100 -1965
<< metal1 >>
rect -3112 1999 -1920 2005
rect -3112 1965 -3100 1999
rect -1932 1965 -1920 1999
rect -3112 1959 -1920 1965
rect -1854 1999 -662 2005
rect -1854 1965 -1842 1999
rect -674 1965 -662 1999
rect -1854 1959 -662 1965
rect -596 1999 596 2005
rect -596 1965 -584 1999
rect 584 1965 596 1999
rect -596 1959 596 1965
rect 662 1999 1854 2005
rect 662 1965 674 1999
rect 1842 1965 1854 1999
rect 662 1959 1854 1965
rect 1920 1999 3112 2005
rect 1920 1965 1932 1999
rect 3100 1965 3112 1999
rect 1920 1959 3112 1965
rect -3168 1915 -3122 1927
rect -3168 1139 -3162 1915
rect -3128 1139 -3122 1915
rect -3168 1127 -3122 1139
rect -1910 1915 -1864 1927
rect -1910 1139 -1904 1915
rect -1870 1139 -1864 1915
rect -1910 1127 -1864 1139
rect -652 1915 -606 1927
rect -652 1139 -646 1915
rect -612 1139 -606 1915
rect -652 1127 -606 1139
rect 606 1915 652 1927
rect 606 1139 612 1915
rect 646 1139 652 1915
rect 606 1127 652 1139
rect 1864 1915 1910 1927
rect 1864 1139 1870 1915
rect 1904 1139 1910 1915
rect 1864 1127 1910 1139
rect 3122 1915 3168 1927
rect 3122 1139 3128 1915
rect 3162 1139 3168 1915
rect 3122 1127 3168 1139
rect -3112 1089 -1920 1095
rect -3112 1055 -3100 1089
rect -1932 1055 -1920 1089
rect -3112 1049 -1920 1055
rect -1854 1089 -662 1095
rect -1854 1055 -1842 1089
rect -674 1055 -662 1089
rect -1854 1049 -662 1055
rect -596 1089 596 1095
rect -596 1055 -584 1089
rect 584 1055 596 1089
rect -596 1049 596 1055
rect 662 1089 1854 1095
rect 662 1055 674 1089
rect 1842 1055 1854 1089
rect 662 1049 1854 1055
rect 1920 1089 3112 1095
rect 1920 1055 1932 1089
rect 3100 1055 3112 1089
rect 1920 1049 3112 1055
rect -3112 981 -1920 987
rect -3112 947 -3100 981
rect -1932 947 -1920 981
rect -3112 941 -1920 947
rect -1854 981 -662 987
rect -1854 947 -1842 981
rect -674 947 -662 981
rect -1854 941 -662 947
rect -596 981 596 987
rect -596 947 -584 981
rect 584 947 596 981
rect -596 941 596 947
rect 662 981 1854 987
rect 662 947 674 981
rect 1842 947 1854 981
rect 662 941 1854 947
rect 1920 981 3112 987
rect 1920 947 1932 981
rect 3100 947 3112 981
rect 1920 941 3112 947
rect -3168 897 -3122 909
rect -3168 121 -3162 897
rect -3128 121 -3122 897
rect -3168 109 -3122 121
rect -1910 897 -1864 909
rect -1910 121 -1904 897
rect -1870 121 -1864 897
rect -1910 109 -1864 121
rect -652 897 -606 909
rect -652 121 -646 897
rect -612 121 -606 897
rect -652 109 -606 121
rect 606 897 652 909
rect 606 121 612 897
rect 646 121 652 897
rect 606 109 652 121
rect 1864 897 1910 909
rect 1864 121 1870 897
rect 1904 121 1910 897
rect 1864 109 1910 121
rect 3122 897 3168 909
rect 3122 121 3128 897
rect 3162 121 3168 897
rect 3122 109 3168 121
rect -3112 71 -1920 77
rect -3112 37 -3100 71
rect -1932 37 -1920 71
rect -3112 31 -1920 37
rect -1854 71 -662 77
rect -1854 37 -1842 71
rect -674 37 -662 71
rect -1854 31 -662 37
rect -596 71 596 77
rect -596 37 -584 71
rect 584 37 596 71
rect -596 31 596 37
rect 662 71 1854 77
rect 662 37 674 71
rect 1842 37 1854 71
rect 662 31 1854 37
rect 1920 71 3112 77
rect 1920 37 1932 71
rect 3100 37 3112 71
rect 1920 31 3112 37
rect -3112 -37 -1920 -31
rect -3112 -71 -3100 -37
rect -1932 -71 -1920 -37
rect -3112 -77 -1920 -71
rect -1854 -37 -662 -31
rect -1854 -71 -1842 -37
rect -674 -71 -662 -37
rect -1854 -77 -662 -71
rect -596 -37 596 -31
rect -596 -71 -584 -37
rect 584 -71 596 -37
rect -596 -77 596 -71
rect 662 -37 1854 -31
rect 662 -71 674 -37
rect 1842 -71 1854 -37
rect 662 -77 1854 -71
rect 1920 -37 3112 -31
rect 1920 -71 1932 -37
rect 3100 -71 3112 -37
rect 1920 -77 3112 -71
rect -3168 -121 -3122 -109
rect -3168 -897 -3162 -121
rect -3128 -897 -3122 -121
rect -3168 -909 -3122 -897
rect -1910 -121 -1864 -109
rect -1910 -897 -1904 -121
rect -1870 -897 -1864 -121
rect -1910 -909 -1864 -897
rect -652 -121 -606 -109
rect -652 -897 -646 -121
rect -612 -897 -606 -121
rect -652 -909 -606 -897
rect 606 -121 652 -109
rect 606 -897 612 -121
rect 646 -897 652 -121
rect 606 -909 652 -897
rect 1864 -121 1910 -109
rect 1864 -897 1870 -121
rect 1904 -897 1910 -121
rect 1864 -909 1910 -897
rect 3122 -121 3168 -109
rect 3122 -897 3128 -121
rect 3162 -897 3168 -121
rect 3122 -909 3168 -897
rect -3112 -947 -1920 -941
rect -3112 -981 -3100 -947
rect -1932 -981 -1920 -947
rect -3112 -987 -1920 -981
rect -1854 -947 -662 -941
rect -1854 -981 -1842 -947
rect -674 -981 -662 -947
rect -1854 -987 -662 -981
rect -596 -947 596 -941
rect -596 -981 -584 -947
rect 584 -981 596 -947
rect -596 -987 596 -981
rect 662 -947 1854 -941
rect 662 -981 674 -947
rect 1842 -981 1854 -947
rect 662 -987 1854 -981
rect 1920 -947 3112 -941
rect 1920 -981 1932 -947
rect 3100 -981 3112 -947
rect 1920 -987 3112 -981
rect -3112 -1055 -1920 -1049
rect -3112 -1089 -3100 -1055
rect -1932 -1089 -1920 -1055
rect -3112 -1095 -1920 -1089
rect -1854 -1055 -662 -1049
rect -1854 -1089 -1842 -1055
rect -674 -1089 -662 -1055
rect -1854 -1095 -662 -1089
rect -596 -1055 596 -1049
rect -596 -1089 -584 -1055
rect 584 -1089 596 -1055
rect -596 -1095 596 -1089
rect 662 -1055 1854 -1049
rect 662 -1089 674 -1055
rect 1842 -1089 1854 -1055
rect 662 -1095 1854 -1089
rect 1920 -1055 3112 -1049
rect 1920 -1089 1932 -1055
rect 3100 -1089 3112 -1055
rect 1920 -1095 3112 -1089
rect -3168 -1139 -3122 -1127
rect -3168 -1915 -3162 -1139
rect -3128 -1915 -3122 -1139
rect -3168 -1927 -3122 -1915
rect -1910 -1139 -1864 -1127
rect -1910 -1915 -1904 -1139
rect -1870 -1915 -1864 -1139
rect -1910 -1927 -1864 -1915
rect -652 -1139 -606 -1127
rect -652 -1915 -646 -1139
rect -612 -1915 -606 -1139
rect -652 -1927 -606 -1915
rect 606 -1139 652 -1127
rect 606 -1915 612 -1139
rect 646 -1915 652 -1139
rect 606 -1927 652 -1915
rect 1864 -1139 1910 -1127
rect 1864 -1915 1870 -1139
rect 1904 -1915 1910 -1139
rect 1864 -1927 1910 -1915
rect 3122 -1139 3168 -1127
rect 3122 -1915 3128 -1139
rect 3162 -1915 3168 -1139
rect 3122 -1927 3168 -1915
rect -3112 -1965 -1920 -1959
rect -3112 -1999 -3100 -1965
rect -1932 -1999 -1920 -1965
rect -3112 -2005 -1920 -1999
rect -1854 -1965 -662 -1959
rect -1854 -1999 -1842 -1965
rect -674 -1999 -662 -1965
rect -1854 -2005 -662 -1999
rect -596 -1965 596 -1959
rect -596 -1999 -584 -1965
rect 584 -1999 596 -1965
rect -596 -2005 596 -1999
rect 662 -1965 1854 -1959
rect 662 -1999 674 -1965
rect 1842 -1999 1854 -1965
rect 662 -2005 1854 -1999
rect 1920 -1965 3112 -1959
rect 1920 -1999 1932 -1965
rect 3100 -1999 3112 -1965
rect 1920 -2005 3112 -1999
<< properties >>
string FIXED_BBOX -3259 -2084 3259 2084
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 6 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
