magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< error_p >>
rect -221 581 -163 587
rect -29 581 29 587
rect 163 581 221 587
rect -221 547 -209 581
rect -29 547 -17 581
rect 163 547 175 581
rect -221 541 -163 547
rect -29 541 29 547
rect 163 541 221 547
rect -125 71 -67 77
rect 67 71 125 77
rect -125 37 -113 71
rect 67 37 79 71
rect -125 31 -67 37
rect 67 31 125 37
rect -125 -37 -67 -31
rect 67 -37 125 -31
rect -125 -71 -113 -37
rect 67 -71 79 -37
rect -125 -77 -67 -71
rect 67 -77 125 -71
rect -221 -547 -163 -541
rect -29 -547 29 -541
rect 163 -547 221 -541
rect -221 -581 -209 -547
rect -29 -581 -17 -547
rect 163 -581 175 -547
rect -221 -587 -163 -581
rect -29 -587 29 -581
rect 163 -587 221 -581
<< pwell >>
rect -407 -719 407 719
<< nmos >>
rect -207 109 -177 509
rect -111 109 -81 509
rect -15 109 15 509
rect 81 109 111 509
rect 177 109 207 509
rect -207 -509 -177 -109
rect -111 -509 -81 -109
rect -15 -509 15 -109
rect 81 -509 111 -109
rect 177 -509 207 -109
<< ndiff >>
rect -269 497 -207 509
rect -269 121 -257 497
rect -223 121 -207 497
rect -269 109 -207 121
rect -177 497 -111 509
rect -177 121 -161 497
rect -127 121 -111 497
rect -177 109 -111 121
rect -81 497 -15 509
rect -81 121 -65 497
rect -31 121 -15 497
rect -81 109 -15 121
rect 15 497 81 509
rect 15 121 31 497
rect 65 121 81 497
rect 15 109 81 121
rect 111 497 177 509
rect 111 121 127 497
rect 161 121 177 497
rect 111 109 177 121
rect 207 497 269 509
rect 207 121 223 497
rect 257 121 269 497
rect 207 109 269 121
rect -269 -121 -207 -109
rect -269 -497 -257 -121
rect -223 -497 -207 -121
rect -269 -509 -207 -497
rect -177 -121 -111 -109
rect -177 -497 -161 -121
rect -127 -497 -111 -121
rect -177 -509 -111 -497
rect -81 -121 -15 -109
rect -81 -497 -65 -121
rect -31 -497 -15 -121
rect -81 -509 -15 -497
rect 15 -121 81 -109
rect 15 -497 31 -121
rect 65 -497 81 -121
rect 15 -509 81 -497
rect 111 -121 177 -109
rect 111 -497 127 -121
rect 161 -497 177 -121
rect 111 -509 177 -497
rect 207 -121 269 -109
rect 207 -497 223 -121
rect 257 -497 269 -121
rect 207 -509 269 -497
<< ndiffc >>
rect -257 121 -223 497
rect -161 121 -127 497
rect -65 121 -31 497
rect 31 121 65 497
rect 127 121 161 497
rect 223 121 257 497
rect -257 -497 -223 -121
rect -161 -497 -127 -121
rect -65 -497 -31 -121
rect 31 -497 65 -121
rect 127 -497 161 -121
rect 223 -497 257 -121
<< psubdiff >>
rect -371 649 -275 683
rect 275 649 371 683
rect -371 587 -337 649
rect 337 587 371 649
rect -371 -649 -337 -587
rect 337 -649 371 -587
rect -371 -683 -275 -649
rect 275 -683 371 -649
<< psubdiffcont >>
rect -275 649 275 683
rect -371 -587 -337 587
rect 337 -587 371 587
rect -275 -683 275 -649
<< poly >>
rect -225 581 -159 597
rect -225 547 -209 581
rect -175 547 -159 581
rect -225 531 -159 547
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -207 509 -177 531
rect -111 509 -81 535
rect -33 531 33 547
rect 159 581 225 597
rect 159 547 175 581
rect 209 547 225 581
rect -15 509 15 531
rect 81 509 111 535
rect 159 531 225 547
rect 177 509 207 531
rect -207 83 -177 109
rect -111 87 -81 109
rect -129 71 -63 87
rect -15 83 15 109
rect 81 87 111 109
rect -129 37 -113 71
rect -79 37 -63 71
rect -129 21 -63 37
rect 63 71 129 87
rect 177 83 207 109
rect 63 37 79 71
rect 113 37 129 71
rect 63 21 129 37
rect -129 -37 -63 -21
rect -129 -71 -113 -37
rect -79 -71 -63 -37
rect -207 -109 -177 -83
rect -129 -87 -63 -71
rect 63 -37 129 -21
rect 63 -71 79 -37
rect 113 -71 129 -37
rect -111 -109 -81 -87
rect -15 -109 15 -83
rect 63 -87 129 -71
rect 81 -109 111 -87
rect 177 -109 207 -83
rect -207 -531 -177 -509
rect -225 -547 -159 -531
rect -111 -535 -81 -509
rect -15 -531 15 -509
rect -225 -581 -209 -547
rect -175 -581 -159 -547
rect -225 -597 -159 -581
rect -33 -547 33 -531
rect 81 -535 111 -509
rect 177 -531 207 -509
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
rect 159 -547 225 -531
rect 159 -581 175 -547
rect 209 -581 225 -547
rect 159 -597 225 -581
<< polycont >>
rect -209 547 -175 581
rect -17 547 17 581
rect 175 547 209 581
rect -113 37 -79 71
rect 79 37 113 71
rect -113 -71 -79 -37
rect 79 -71 113 -37
rect -209 -581 -175 -547
rect -17 -581 17 -547
rect 175 -581 209 -547
<< locali >>
rect -371 649 -275 683
rect 275 649 371 683
rect -371 587 -337 649
rect 337 587 371 649
rect -225 547 -209 581
rect -175 547 -159 581
rect -33 547 -17 581
rect 17 547 33 581
rect 159 547 175 581
rect 209 547 225 581
rect -257 497 -223 513
rect -257 105 -223 121
rect -161 497 -127 513
rect -161 105 -127 121
rect -65 497 -31 513
rect -65 105 -31 121
rect 31 497 65 513
rect 31 105 65 121
rect 127 497 161 513
rect 127 105 161 121
rect 223 497 257 513
rect 223 105 257 121
rect -129 37 -113 71
rect -79 37 -63 71
rect 63 37 79 71
rect 113 37 129 71
rect -129 -71 -113 -37
rect -79 -71 -63 -37
rect 63 -71 79 -37
rect 113 -71 129 -37
rect -257 -121 -223 -105
rect -257 -513 -223 -497
rect -161 -121 -127 -105
rect -161 -513 -127 -497
rect -65 -121 -31 -105
rect -65 -513 -31 -497
rect 31 -121 65 -105
rect 31 -513 65 -497
rect 127 -121 161 -105
rect 127 -513 161 -497
rect 223 -121 257 -105
rect 223 -513 257 -497
rect -225 -581 -209 -547
rect -175 -581 -159 -547
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect 159 -581 175 -547
rect 209 -581 225 -547
rect -371 -649 -337 -587
rect 337 -649 371 -587
rect -371 -683 -275 -649
rect 275 -683 371 -649
<< viali >>
rect -209 547 -175 581
rect -17 547 17 581
rect 175 547 209 581
rect -257 121 -223 497
rect -161 121 -127 497
rect -65 121 -31 497
rect 31 121 65 497
rect 127 121 161 497
rect 223 121 257 497
rect -113 37 -79 71
rect 79 37 113 71
rect -113 -71 -79 -37
rect 79 -71 113 -37
rect -257 -497 -223 -121
rect -161 -497 -127 -121
rect -65 -497 -31 -121
rect 31 -497 65 -121
rect 127 -497 161 -121
rect 223 -497 257 -121
rect -209 -581 -175 -547
rect -17 -581 17 -547
rect 175 -581 209 -547
<< metal1 >>
rect -221 581 -163 587
rect -221 547 -209 581
rect -175 547 -163 581
rect -221 541 -163 547
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect 163 581 221 587
rect 163 547 175 581
rect 209 547 221 581
rect 163 541 221 547
rect -263 497 -217 509
rect -263 121 -257 497
rect -223 121 -217 497
rect -263 109 -217 121
rect -167 497 -121 509
rect -167 121 -161 497
rect -127 121 -121 497
rect -167 109 -121 121
rect -71 497 -25 509
rect -71 121 -65 497
rect -31 121 -25 497
rect -71 109 -25 121
rect 25 497 71 509
rect 25 121 31 497
rect 65 121 71 497
rect 25 109 71 121
rect 121 497 167 509
rect 121 121 127 497
rect 161 121 167 497
rect 121 109 167 121
rect 217 497 263 509
rect 217 121 223 497
rect 257 121 263 497
rect 217 109 263 121
rect -125 71 -67 77
rect -125 37 -113 71
rect -79 37 -67 71
rect -125 31 -67 37
rect 67 71 125 77
rect 67 37 79 71
rect 113 37 125 71
rect 67 31 125 37
rect -125 -37 -67 -31
rect -125 -71 -113 -37
rect -79 -71 -67 -37
rect -125 -77 -67 -71
rect 67 -37 125 -31
rect 67 -71 79 -37
rect 113 -71 125 -37
rect 67 -77 125 -71
rect -263 -121 -217 -109
rect -263 -497 -257 -121
rect -223 -497 -217 -121
rect -263 -509 -217 -497
rect -167 -121 -121 -109
rect -167 -497 -161 -121
rect -127 -497 -121 -121
rect -167 -509 -121 -497
rect -71 -121 -25 -109
rect -71 -497 -65 -121
rect -31 -497 -25 -121
rect -71 -509 -25 -497
rect 25 -121 71 -109
rect 25 -497 31 -121
rect 65 -497 71 -121
rect 25 -509 71 -497
rect 121 -121 167 -109
rect 121 -497 127 -121
rect 161 -497 167 -121
rect 121 -509 167 -497
rect 217 -121 263 -109
rect 217 -497 223 -121
rect 257 -497 263 -121
rect 217 -509 263 -497
rect -221 -547 -163 -541
rect -221 -581 -209 -547
rect -175 -581 -163 -547
rect -221 -587 -163 -581
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
rect 163 -547 221 -541
rect 163 -581 175 -547
rect 209 -581 221 -547
rect 163 -587 221 -581
<< properties >>
string FIXED_BBOX -354 -666 354 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
