magic
tech sky130A
magscale 1 2
timestamp 1645789405
<< pwell >>
rect -941 -810 941 810
<< nmos >>
rect -745 -600 -545 600
rect -487 -600 -287 600
rect -229 -600 -29 600
rect 29 -600 229 600
rect 287 -600 487 600
rect 545 -600 745 600
<< ndiff >>
rect -803 588 -745 600
rect -803 -588 -791 588
rect -757 -588 -745 588
rect -803 -600 -745 -588
rect -545 588 -487 600
rect -545 -588 -533 588
rect -499 -588 -487 588
rect -545 -600 -487 -588
rect -287 588 -229 600
rect -287 -588 -275 588
rect -241 -588 -229 588
rect -287 -600 -229 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 229 588 287 600
rect 229 -588 241 588
rect 275 -588 287 588
rect 229 -600 287 -588
rect 487 588 545 600
rect 487 -588 499 588
rect 533 -588 545 588
rect 487 -600 545 -588
rect 745 588 803 600
rect 745 -588 757 588
rect 791 -588 803 588
rect 745 -600 803 -588
<< ndiffc >>
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
<< psubdiff >>
rect -905 740 -809 774
rect 809 740 905 774
rect -905 678 -871 740
rect 871 678 905 740
rect -905 -740 -871 -678
rect 871 -740 905 -678
rect -905 -774 -809 -740
rect 809 -774 905 -740
<< psubdiffcont >>
rect -809 740 809 774
rect -905 -678 -871 678
rect 871 -678 905 678
rect -809 -774 809 -740
<< poly >>
rect -745 672 -545 688
rect -745 638 -729 672
rect -561 638 -545 672
rect -745 600 -545 638
rect -487 672 -287 688
rect -487 638 -471 672
rect -303 638 -287 672
rect -487 600 -287 638
rect -229 672 -29 688
rect -229 638 -213 672
rect -45 638 -29 672
rect -229 600 -29 638
rect 29 672 229 688
rect 29 638 45 672
rect 213 638 229 672
rect 29 600 229 638
rect 287 672 487 688
rect 287 638 303 672
rect 471 638 487 672
rect 287 600 487 638
rect 545 672 745 688
rect 545 638 561 672
rect 729 638 745 672
rect 545 600 745 638
rect -745 -638 -545 -600
rect -745 -672 -729 -638
rect -561 -672 -545 -638
rect -745 -688 -545 -672
rect -487 -638 -287 -600
rect -487 -672 -471 -638
rect -303 -672 -287 -638
rect -487 -688 -287 -672
rect -229 -638 -29 -600
rect -229 -672 -213 -638
rect -45 -672 -29 -638
rect -229 -688 -29 -672
rect 29 -638 229 -600
rect 29 -672 45 -638
rect 213 -672 229 -638
rect 29 -688 229 -672
rect 287 -638 487 -600
rect 287 -672 303 -638
rect 471 -672 487 -638
rect 287 -688 487 -672
rect 545 -638 745 -600
rect 545 -672 561 -638
rect 729 -672 745 -638
rect 545 -688 745 -672
<< polycont >>
rect -729 638 -561 672
rect -471 638 -303 672
rect -213 638 -45 672
rect 45 638 213 672
rect 303 638 471 672
rect 561 638 729 672
rect -729 -672 -561 -638
rect -471 -672 -303 -638
rect -213 -672 -45 -638
rect 45 -672 213 -638
rect 303 -672 471 -638
rect 561 -672 729 -638
<< locali >>
rect -905 740 -809 774
rect 809 740 905 774
rect -905 678 -871 740
rect 871 678 905 740
rect -745 638 -729 672
rect -561 638 -545 672
rect -487 638 -471 672
rect -303 638 -287 672
rect -229 638 -213 672
rect -45 638 -29 672
rect 29 638 45 672
rect 213 638 229 672
rect 287 638 303 672
rect 471 638 487 672
rect 545 638 561 672
rect 729 638 745 672
rect -791 588 -757 604
rect -791 -604 -757 -588
rect -533 588 -499 604
rect -533 -604 -499 -588
rect -275 588 -241 604
rect -275 -604 -241 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 241 588 275 604
rect 241 -604 275 -588
rect 499 588 533 604
rect 499 -604 533 -588
rect 757 588 791 604
rect 757 -604 791 -588
rect -745 -672 -729 -638
rect -561 -672 -545 -638
rect -487 -672 -471 -638
rect -303 -672 -287 -638
rect -229 -672 -213 -638
rect -45 -672 -29 -638
rect 29 -672 45 -638
rect 213 -672 229 -638
rect 287 -672 303 -638
rect 471 -672 487 -638
rect 545 -672 561 -638
rect 729 -672 745 -638
rect -905 -740 -871 -678
rect 871 -740 905 -678
rect -905 -774 -809 -740
rect 809 -774 905 -740
<< viali >>
rect -729 638 -561 672
rect -471 638 -303 672
rect -213 638 -45 672
rect 45 638 213 672
rect 303 638 471 672
rect 561 638 729 672
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect -729 -672 -561 -638
rect -471 -672 -303 -638
rect -213 -672 -45 -638
rect 45 -672 213 -638
rect 303 -672 471 -638
rect 561 -672 729 -638
<< metal1 >>
rect -741 672 -549 678
rect -741 638 -729 672
rect -561 638 -549 672
rect -741 632 -549 638
rect -483 672 -291 678
rect -483 638 -471 672
rect -303 638 -291 672
rect -483 632 -291 638
rect -225 672 -33 678
rect -225 638 -213 672
rect -45 638 -33 672
rect -225 632 -33 638
rect 33 672 225 678
rect 33 638 45 672
rect 213 638 225 672
rect 33 632 225 638
rect 291 672 483 678
rect 291 638 303 672
rect 471 638 483 672
rect 291 632 483 638
rect 549 672 741 678
rect 549 638 561 672
rect 729 638 741 672
rect 549 632 741 638
rect -797 588 -751 600
rect -797 -588 -791 588
rect -757 -588 -751 588
rect -797 -600 -751 -588
rect -539 588 -493 600
rect -539 -588 -533 588
rect -499 -588 -493 588
rect -539 -600 -493 -588
rect -281 588 -235 600
rect -281 -588 -275 588
rect -241 -588 -235 588
rect -281 -600 -235 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 235 588 281 600
rect 235 -588 241 588
rect 275 -588 281 588
rect 235 -600 281 -588
rect 493 588 539 600
rect 493 -588 499 588
rect 533 -588 539 588
rect 493 -600 539 -588
rect 751 588 797 600
rect 751 -588 757 588
rect 791 -588 797 588
rect 751 -600 797 -588
rect -741 -638 -549 -632
rect -741 -672 -729 -638
rect -561 -672 -549 -638
rect -741 -678 -549 -672
rect -483 -638 -291 -632
rect -483 -672 -471 -638
rect -303 -672 -291 -638
rect -483 -678 -291 -672
rect -225 -638 -33 -632
rect -225 -672 -213 -638
rect -45 -672 -33 -638
rect -225 -678 -33 -672
rect 33 -638 225 -632
rect 33 -672 45 -638
rect 213 -672 225 -638
rect 33 -678 225 -672
rect 291 -638 483 -632
rect 291 -672 303 -638
rect 471 -672 483 -638
rect 291 -678 483 -672
rect 549 -638 741 -632
rect 549 -672 561 -638
rect 729 -672 741 -638
rect 549 -678 741 -672
<< properties >>
string FIXED_BBOX -888 -757 888 757
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
