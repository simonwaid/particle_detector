magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< locali >>
rect -10 70 100 630
rect 630 70 740 630
rect -20 -20 750 70
<< metal1 >>
rect 130 670 600 720
rect 70 460 80 630
rect 140 460 150 630
rect 190 190 240 670
rect 580 460 590 630
rect 650 460 660 630
rect 320 230 330 410
rect 400 230 410 410
rect 130 140 600 190
rect 190 -100 240 140
rect -50 -150 1110 -100
rect -50 -630 10 -150
rect 60 -360 70 -190
rect 130 -360 140 -190
rect 320 -360 330 -190
rect 390 -360 400 -190
rect 580 -360 590 -190
rect 650 -360 660 -190
rect 830 -360 840 -190
rect 900 -360 910 -190
rect 1090 -360 1100 -190
rect 1160 -360 1170 -190
rect 190 -590 200 -420
rect 260 -590 270 -420
rect 450 -590 460 -420
rect 520 -590 530 -420
rect 710 -590 720 -420
rect 780 -590 790 -420
rect 960 -590 970 -420
rect 1030 -590 1040 -420
rect -50 -680 1110 -630
<< via1 >>
rect 80 460 140 630
rect 590 460 650 630
rect 330 230 400 410
rect 70 -360 130 -190
rect 330 -360 390 -190
rect 590 -360 650 -190
rect 840 -360 900 -190
rect 1100 -360 1160 -190
rect 200 -590 260 -420
rect 460 -590 520 -420
rect 720 -590 780 -420
rect 970 -590 1030 -420
<< metal2 >>
rect 80 630 650 640
rect 140 470 590 630
rect 80 450 140 460
rect 590 450 650 460
rect 330 410 400 420
rect 290 230 330 330
rect 400 230 440 330
rect 70 -190 130 -180
rect 290 -190 440 230
rect 590 -190 650 -180
rect 840 -190 900 -180
rect 1100 -190 1160 -180
rect 130 -340 330 -190
rect 70 -370 130 -360
rect 390 -340 590 -190
rect 330 -370 390 -360
rect 650 -340 840 -190
rect 590 -370 650 -360
rect 900 -340 1100 -190
rect 840 -370 900 -360
rect 1100 -370 1160 -360
rect 200 -420 260 -410
rect 460 -420 520 -410
rect 260 -590 460 -440
rect 720 -420 780 -410
rect 520 -590 720 -440
rect 970 -420 1030 -410
rect 780 -590 970 -440
rect 200 -600 260 -590
rect 460 -600 520 -590
rect 720 -600 780 -590
rect 970 -600 1030 -590
use sky130_fd_pr__pfet_01v8_lvt_4LMUGG  sky130_fd_pr__pfet_01v8_lvt_4LMUGG_0
timestamp 1654768133
transform 1 0 619 0 1 -391
box -679 -419 679 419
use sky130_fd_pr__pfet_01v8_lvt_LKHJAY  sky130_fd_pr__pfet_01v8_lvt_LKHJAY_0
timestamp 1654768133
transform 1 0 365 0 1 429
box -425 -419 425 419
<< end >>
