VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mirror_n
  CLASS BLOCK ;
  FOREIGN mirror_n ;
  ORIGIN 0.150 0.150 ;
  SIZE 4.250 BY 17.400 ;
  OBS
      LAYER pwell ;
        RECT -0.150 13.220 2.500 17.250 ;
        RECT -0.150 -0.150 4.100 13.220 ;
      LAYER li1 ;
        RECT -0.150 -0.150 4.100 17.250 ;
      LAYER met1 ;
        RECT 0.500 0.450 3.450 16.700 ;
      LAYER met2 ;
        RECT 0.050 -0.150 3.850 16.250 ;
  END
END mirror_n
MACRO mirror_p
  CLASS BLOCK ;
  FOREIGN mirror_p ;
  ORIGIN 1.600 9.400 ;
  SIZE 6.850 BY 17.900 ;
  OBS
      LAYER nwell ;
        RECT -1.600 4.330 2.030 8.490 ;
        RECT -1.600 -9.400 5.230 4.330 ;
      LAYER li1 ;
        RECT -1.600 -9.400 5.250 8.500 ;
      LAYER met1 ;
        RECT -0.950 -8.750 4.580 7.950 ;
      LAYER met2 ;
        RECT -1.200 -8.400 4.800 7.450 ;
      LAYER met3 ;
        RECT -1.250 -9.400 4.850 6.275 ;
  END
END mirror_p
MACRO sky130_fd_pr__cap_mim_m3_2_LJ5JLG
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_mim_m3_2_LJ5JLG ;
  ORIGIN 16.755 15.500 ;
  SIZE 31.000 BY 31.000 ;
  OBS
      LAYER met4 ;
        RECT -16.755 -15.500 16.755 15.500 ;
      LAYER met5 ;
        RECT -16.175 -15.500 14.245 15.500 ;
        RECT 15.265 -15.505 16.865 15.505 ;
  END
END sky130_fd_pr__cap_mim_m3_2_LJ5JLG
MACRO cmirror_channel
  CLASS BLOCK ;
  FOREIGN cmirror_channel ;
  ORIGIN 0.300 55.500 ;
  SIZE 99.510 BY 76.120 ;
  OBS
      LAYER li1 ;
        RECT 3.300 -19.150 96.850 16.650 ;
      LAYER met1 ;
        RECT -0.300 -21.550 96.200 16.000 ;
      LAYER met2 ;
        RECT -0.250 -21.600 96.450 15.650 ;
      LAYER met3 ;
        RECT -0.300 -21.575 96.850 20.600 ;
      LAYER met4 ;
        RECT -0.255 -55.390 99.205 20.505 ;
      LAYER met5 ;
        RECT 2.750 -55.500 99.210 20.620 ;
  END
END cmirror_channel
END LIBRARY

