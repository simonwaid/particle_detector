* SPICE3 file created from outd_flat.ext - technology: sky130A

X0 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X7 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X10 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X14 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X15 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X19 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X21 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X22 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X23 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X24 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X26 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X28 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X29 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X33 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X36 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X38 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X39 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X40 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X41 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X42 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X43 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X44 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X45 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X46 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X47 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X48 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X51 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X52 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X53 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X54 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X55 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X56 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X57 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X58 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X59 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X61 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X62 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X63 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X64 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X65 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X66 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X67 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X69 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X70 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X71 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X72 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X75 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X76 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X77 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X80 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X82 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X83 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X84 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X85 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X86 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X87 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X90 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X92 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X93 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X94 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X95 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X98 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X99 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X100 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X101 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X102 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X104 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X105 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X106 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X107 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X108 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X109 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X110 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X111 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X112 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X113 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X114 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X115 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X116 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X117 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X118 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X119 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X120 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X121 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X122 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X123 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X124 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X125 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X126 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X127 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X128 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X129 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X130 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X131 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X132 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X133 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X134 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X135 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X136 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X137 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X138 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X139 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X140 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X141 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X142 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X143 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X145 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X146 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X147 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X148 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X149 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X150 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X151 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X152 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X153 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X154 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X155 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X156 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X157 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X158 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X159 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X160 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X161 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X162 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X163 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X164 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X165 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X166 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X167 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X168 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X169 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X170 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X171 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X172 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X173 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X174 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X175 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X176 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X177 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X178 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X179 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X180 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X181 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X182 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X183 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X184 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X185 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X186 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X187 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X188 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X189 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X190 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X191 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X192 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X193 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X194 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X195 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X196 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X197 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X198 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X199 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X200 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X201 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X202 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X203 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X204 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X205 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X206 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X207 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X208 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X209 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X210 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X211 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X212 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X213 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X214 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X215 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X216 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X217 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X218 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X219 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X220 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X221 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X222 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X223 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X224 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X225 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X226 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X227 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X228 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X229 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X230 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X231 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X232 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X233 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X234 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X235 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X236 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X237 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X238 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X239 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X240 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X241 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X242 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X243 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X244 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X245 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X246 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X247 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X248 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X249 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X250 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X251 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X252 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X253 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X254 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X255 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X256 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X257 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X258 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X259 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X261 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X262 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X263 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X264 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X265 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X266 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X267 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X268 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X269 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X273 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X274 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X275 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X276 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X277 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X279 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X280 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X281 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X283 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X284 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X285 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X286 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X287 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X288 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X289 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X290 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X291 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X292 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X293 V_da2_N VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X294 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X295 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X296 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X297 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X298 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X299 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X300 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X301 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X302 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X303 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X304 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X305 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X306 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X307 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X308 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X309 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X310 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X311 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X312 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X313 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X314 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X315 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X316 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X317 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X318 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X319 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X320 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X321 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X322 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X323 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X324 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X325 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X326 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X327 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X328 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X329 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X330 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X331 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X332 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X333 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X334 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X335 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X336 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X337 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X338 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X339 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X340 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X341 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X342 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X343 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X344 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X345 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X346 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X347 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X348 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X349 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X350 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X351 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X352 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X353 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X354 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X355 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X356 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X357 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X358 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X359 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X360 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X361 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X362 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X363 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X364 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X365 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X366 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X367 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X368 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X369 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X370 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X371 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X372 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X373 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X374 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X375 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X376 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X377 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X378 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X379 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X380 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X381 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X382 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X383 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X384 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X385 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X386 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X387 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X388 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X389 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X390 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X391 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X392 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X393 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X394 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X395 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X396 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X397 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X398 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X399 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X400 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X401 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X402 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X403 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X404 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X405 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X406 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X407 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X408 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X409 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X410 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X411 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X412 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X413 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X414 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X415 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X416 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X417 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X418 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X419 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X420 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X421 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X422 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X423 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X424 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X425 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X426 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X427 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X428 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X429 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X430 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X431 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X432 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X433 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X434 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X435 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X436 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X437 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X438 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X439 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X440 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X441 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X442 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X443 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X444 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X445 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X446 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X447 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X448 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X449 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X450 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X451 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X452 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X453 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X454 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X455 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X456 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X457 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X458 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X459 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X460 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X461 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X462 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X463 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X464 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X465 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X466 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X467 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X468 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X469 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X470 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X471 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X472 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X473 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X474 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X475 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X476 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X477 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X478 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X479 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X480 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X481 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X482 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X483 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X484 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X485 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X486 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X487 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X488 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X489 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X490 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X491 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X492 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X493 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X494 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X495 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X496 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X497 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X498 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X499 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X500 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X501 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X502 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X503 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X504 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X505 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X506 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X507 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X508 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X509 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X510 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X511 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X512 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X513 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X514 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X515 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X516 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X517 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X519 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X520 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X521 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X522 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X523 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X524 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X525 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X526 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X527 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X528 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X529 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X530 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X531 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X532 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X533 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X534 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X535 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X536 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X537 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X538 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X540 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X541 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X542 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X543 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X544 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X545 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X546 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X547 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X548 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X549 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X550 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X551 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X552 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X553 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X554 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X555 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X556 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X557 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X558 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X559 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X560 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X561 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X562 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X563 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X564 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X565 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X566 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X567 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X568 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X569 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X570 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X571 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X572 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X573 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X574 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X575 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X576 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X577 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X578 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X579 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X580 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X581 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X582 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X583 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X584 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X585 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X586 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X587 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X588 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X589 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X590 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X591 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X592 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X593 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X594 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X595 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X596 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X597 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X598 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X599 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X600 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X601 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X602 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X603 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X604 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X605 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X606 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X607 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X608 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X609 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X610 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X611 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X612 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X613 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X614 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X615 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X616 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X617 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X618 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X619 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X620 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X621 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X622 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X623 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X624 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X625 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X626 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X627 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X628 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X629 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X630 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X631 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X632 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X633 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X634 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X635 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X636 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X637 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X638 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X639 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X640 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X641 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X642 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X643 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X644 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X645 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X646 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X647 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X648 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X649 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X650 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X651 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X652 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X653 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X654 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X655 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X656 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X657 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X658 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X659 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X660 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X661 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X662 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X663 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X664 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X665 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X666 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X667 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X668 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X669 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X670 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X671 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X672 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X673 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X674 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X675 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X676 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X677 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X678 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X679 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X680 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X681 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X682 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X683 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X684 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X685 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X686 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X687 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X688 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X689 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X690 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X691 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X692 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X693 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X694 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X695 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X696 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X697 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X698 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X699 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X700 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X701 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X702 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X703 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X704 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X705 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X706 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X707 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X708 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X709 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X710 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X711 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X712 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X713 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X714 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X715 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X716 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X717 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X718 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X719 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X720 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X721 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X722 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X723 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X724 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X725 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X726 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X727 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X728 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X729 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X730 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X731 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X732 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X733 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X734 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X735 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X736 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X737 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X738 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X739 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X740 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X741 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X742 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X743 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X744 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X745 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X746 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X747 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X748 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X749 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X750 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X751 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X752 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X753 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X754 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X755 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X756 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X757 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X758 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X759 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X760 V_da2_P VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X761 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X762 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X763 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X764 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X765 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X766 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X767 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X768 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X769 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X770 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X771 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X772 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X773 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X774 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X775 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X776 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X777 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X778 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X779 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X780 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X781 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X782 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X783 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X784 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X785 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X786 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X787 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X788 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X789 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X790 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X791 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X792 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X793 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X794 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X795 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X796 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X797 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X798 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X799 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X800 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X801 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X802 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X803 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X804 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X805 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X806 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X807 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X808 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X809 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X810 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X811 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X812 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X813 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X814 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X815 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X816 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X817 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X818 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X819 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X820 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X821 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X822 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X823 VP V_da2_N outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X824 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X825 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X826 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X827 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X828 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X829 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X830 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X831 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X832 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X833 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X834 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X835 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X836 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X837 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X838 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X839 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X840 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X841 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X842 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X843 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X844 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X845 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X846 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X847 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X848 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X849 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X850 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X851 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X852 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X853 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X854 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X855 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X856 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X857 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X858 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X859 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X860 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X861 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X862 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X863 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X864 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X865 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X866 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X867 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X868 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X869 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X870 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X871 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X872 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X873 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X874 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X875 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X876 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X877 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X878 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X879 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X880 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X881 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X882 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X883 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X884 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X885 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X886 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X887 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X888 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X889 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X890 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X891 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X892 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X893 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X894 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X895 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X896 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X897 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X898 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X899 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X900 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X901 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X902 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X903 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X904 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X905 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X906 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X907 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X908 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X909 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X910 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X911 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X912 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X913 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X914 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X915 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X916 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X917 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X918 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X919 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X920 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X921 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X922 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X923 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X924 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X925 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X926 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X927 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X928 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X929 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X930 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X931 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X932 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X933 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X934 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X935 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X936 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X937 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X938 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X939 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X940 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X941 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X942 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X943 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X944 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X945 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X946 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X947 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X948 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X949 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X950 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X951 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X952 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X953 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X954 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X955 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X956 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X957 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X958 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X959 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X960 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X961 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X962 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X963 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X964 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X965 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X966 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X967 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X968 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X969 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X970 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X971 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X972 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X973 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X974 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X975 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X976 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X977 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X978 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X979 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X980 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X981 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X982 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X983 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X984 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X985 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X986 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X987 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X988 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X989 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X990 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X991 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X992 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X993 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X994 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X995 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X996 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X997 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X998 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X999 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1000 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1001 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1002 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1003 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1004 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1005 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1006 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1007 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1008 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1009 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1010 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1011 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1012 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1013 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1014 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1015 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1016 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1017 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1018 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1019 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1020 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1021 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1022 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1023 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1024 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1025 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1026 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1027 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1028 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1029 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1030 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1031 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1032 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1033 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1034 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1035 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1036 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1037 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1038 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1039 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1040 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1041 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1042 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1043 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1044 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1045 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1046 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1047 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1048 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1049 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1050 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1051 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1052 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1053 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1054 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1055 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1056 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1057 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1058 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1059 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1060 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1061 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1062 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1063 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1064 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1065 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1066 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1067 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1068 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1069 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1070 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1071 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1072 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1073 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1074 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1075 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1076 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1077 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1078 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1079 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1080 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1081 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1082 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1083 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1084 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1085 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1086 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1087 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1088 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1089 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1090 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1091 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1092 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1093 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1094 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1095 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1096 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1097 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1098 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1099 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1100 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1101 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1102 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1103 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1104 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1105 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1106 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1107 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1108 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1109 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1110 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1111 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1112 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1113 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1114 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1115 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1116 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1117 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1118 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1119 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1120 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1121 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1122 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1123 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1124 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1125 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1126 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1127 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1128 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1129 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1130 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1131 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1132 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1133 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1134 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1135 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1136 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1137 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1138 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1139 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1140 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1141 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1142 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1143 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1144 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1145 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1146 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1147 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1148 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1149 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1150 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1151 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1152 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1153 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1154 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1155 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1156 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1157 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1158 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1159 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1160 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1161 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1162 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1163 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1164 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1165 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1166 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1167 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1168 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1169 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1170 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1171 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1172 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1173 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1174 V_da2_P VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1175 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1176 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1177 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1178 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1179 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1180 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1181 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1182 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1183 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1184 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1185 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1186 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1187 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1188 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1189 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1190 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1191 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1192 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1193 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1194 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1195 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1196 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1197 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1198 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1199 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1200 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1201 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1202 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1203 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1204 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1205 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1206 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1207 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1208 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1209 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1210 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1211 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1212 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1213 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1214 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1215 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1216 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1217 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1218 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1219 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1220 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1221 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1222 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1223 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1224 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1225 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1226 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1227 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1228 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1229 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1230 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1231 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1232 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1233 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1234 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1235 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1236 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1237 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1238 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1239 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1240 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1241 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1242 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1243 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1244 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1245 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1246 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1247 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1248 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1249 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1250 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1251 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1252 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1253 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1254 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1255 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1256 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1257 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1258 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1259 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1260 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1261 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1262 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1263 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1264 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1265 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1266 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1267 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1268 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1269 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1270 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1271 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1272 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1273 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1274 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1275 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1276 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1277 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1278 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1279 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1280 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1281 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1282 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1283 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1284 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1285 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1286 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1287 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1288 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1289 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1290 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1291 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1292 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1293 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1294 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1295 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1296 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1297 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1298 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1299 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1300 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1301 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1302 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1303 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1304 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1305 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1306 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1307 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1308 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1309 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1310 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1311 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1312 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1313 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1314 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1315 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1316 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1317 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1318 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1319 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1320 V_da2_N VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1321 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1322 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1323 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1324 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1325 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1326 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1327 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1328 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1329 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1330 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1331 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1332 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1333 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1334 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1335 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1336 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1337 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1338 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1339 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1340 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1341 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1342 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1343 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1344 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1345 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1346 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1347 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1348 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1349 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1350 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1351 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1352 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1353 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1354 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1355 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1356 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1357 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1358 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1359 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1360 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1361 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1362 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1363 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1364 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1365 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1366 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1367 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1368 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1369 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1370 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1371 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1372 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1373 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1374 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1375 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1376 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1377 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1378 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1379 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1380 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1381 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1382 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1383 V_da1_N VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X1384 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1385 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1386 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1387 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1388 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1389 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1390 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1391 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1392 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1393 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1394 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1395 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1396 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1397 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1398 V_da1_P VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X1399 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1400 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1401 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1402 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1403 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1404 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1405 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1406 V_da1_N VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X1407 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1408 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1409 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1410 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1411 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1412 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1413 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1414 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1415 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1416 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1417 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1418 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1419 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1420 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1421 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1422 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1423 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1424 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1425 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1426 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1427 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1428 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1429 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1430 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1431 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1432 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1433 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1434 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1435 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1436 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1437 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1438 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1439 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1440 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1441 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1442 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1443 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1444 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1445 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1446 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1447 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1448 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1449 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1450 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1451 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1452 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1453 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1454 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1455 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1456 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1457 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1458 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1459 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1460 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1461 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1462 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1463 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1464 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1465 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1466 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1467 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1468 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1469 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1470 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1471 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1472 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1473 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1474 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1475 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1476 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1477 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1478 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1479 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1480 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1481 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1482 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1483 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1484 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1485 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1486 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1487 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1488 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1489 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1490 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1491 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1492 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1493 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1494 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1495 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1496 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1497 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1498 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1499 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1500 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1501 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1502 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1503 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1504 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1505 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1506 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1507 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1508 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1509 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1510 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1511 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1512 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1513 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1514 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1515 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1516 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1517 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1518 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1519 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1520 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1521 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1522 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1523 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1524 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1525 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1526 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1527 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1528 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1529 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1530 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1531 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1532 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1533 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1534 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1535 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1536 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1537 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1538 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1539 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1540 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1541 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1542 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1543 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1544 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1545 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1546 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1547 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1548 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1549 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1550 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1551 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1552 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1553 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1554 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1555 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1556 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1557 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1558 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1559 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1560 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1561 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1562 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1563 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1564 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1565 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1566 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1567 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1568 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1569 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1570 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1571 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1572 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1573 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1574 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1575 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1576 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1577 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1578 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1579 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1580 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1581 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1582 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1583 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1584 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1585 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1586 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1587 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1588 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1589 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1590 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1591 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1592 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1593 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1594 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1595 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1596 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1597 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1598 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1599 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1600 V_da1_P VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X1601 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1602 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1603 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1604 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1605 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1606 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1607 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1608 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1609 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1610 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1611 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1612 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1613 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1614 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1615 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19882_7120# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1616 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1617 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1618 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1619 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1620 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1621 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1622 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1623 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1624 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1625 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1626 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1627 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1628 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1629 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1630 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1631 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1632 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1633 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1634 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1635 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1636 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1637 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1638 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1639 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1640 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1641 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1642 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1643 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1644 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1645 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1646 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1647 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1648 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1649 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1650 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1651 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1652 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1653 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1654 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1655 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1656 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1657 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1658 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1659 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1660 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1661 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1662 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1663 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1664 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1665 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1666 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1667 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1668 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1669 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1670 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1671 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1672 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1673 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1674 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1675 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1676 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1677 a_n19882_7120# I_Bias I_Bias outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1678 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1679 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1680 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1681 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1682 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1683 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1684 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1685 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1686 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1687 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1688 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1689 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1690 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1691 VP V_da2_P outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1692 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1693 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1694 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1695 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1696 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1697 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1698 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1699 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1700 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1701 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1702 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1703 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1704 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1705 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1706 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1707 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1708 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1709 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1710 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1711 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1712 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1713 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1714 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1715 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1716 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1717 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1718 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1719 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1720 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1721 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1722 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1723 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1724 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1725 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1726 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1727 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1728 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1729 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1730 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1731 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1732 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1733 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1734 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1735 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1736 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1737 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1738 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1739 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1740 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1741 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1742 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1743 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1744 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1745 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1746 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1747 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1748 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1749 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1750 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1751 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1752 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1753 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1754 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1755 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1756 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1757 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1758 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1759 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1760 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1761 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1762 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1763 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1764 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1765 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1766 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1767 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1768 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1769 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1770 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1771 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1772 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1773 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1774 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1775 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1776 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1777 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1778 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1779 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1780 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1781 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1782 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1783 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1784 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1785 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1786 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1787 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1788 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1789 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1790 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1791 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1792 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1793 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1794 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1795 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1796 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1797 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1798 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1799 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1800 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1801 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1802 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1803 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1804 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1805 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1806 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1807 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1808 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1809 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1810 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1811 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1812 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1813 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1814 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1815 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1816 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1817 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1818 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1819 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1820 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1821 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1822 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1823 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1824 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1825 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1826 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1827 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1828 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1829 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1830 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1831 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1832 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1833 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1834 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1835 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1836 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1837 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1838 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1839 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1840 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1841 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1842 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1843 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1844 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1845 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1846 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1847 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1848 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1849 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1850 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1851 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1852 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1853 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1854 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1855 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1856 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1857 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1858 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1859 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1860 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1861 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1862 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1863 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1864 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1865 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1866 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1867 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1868 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1869 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1870 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1871 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1872 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1873 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1874 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1875 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1876 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1877 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1878 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1879 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1880 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1881 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1882 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1883 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1884 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1885 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1886 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1887 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1888 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1889 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1890 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1891 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1892 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1893 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1894 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1895 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1896 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1897 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1898 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1899 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1900 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1901 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1902 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1903 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1904 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1905 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1906 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1907 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1908 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1909 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1910 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1911 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1912 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1913 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1914 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1915 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1916 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1917 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1918 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1919 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1920 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1921 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1922 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1923 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1924 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1925 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1926 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1927 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1928 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1929 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1930 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1931 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1932 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1933 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1934 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1935 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1936 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1937 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1938 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1939 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1940 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1941 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1942 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1943 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1944 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1945 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1946 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1947 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1948 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1949 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1950 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1951 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1952 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1953 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1954 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1955 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1956 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1957 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1958 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1959 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1960 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1961 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1962 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1963 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1964 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1965 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X1966 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1967 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1968 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1969 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1970 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1971 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1972 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1973 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1974 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1975 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1976 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1977 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1978 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1979 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1980 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1981 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1982 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1983 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1984 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1985 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1986 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1987 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1988 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1989 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1990 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1991 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1992 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1993 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1994 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1995 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1996 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1997 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1998 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1999 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2000 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2001 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2002 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2003 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2004 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2005 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2006 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2007 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2008 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2009 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2010 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2011 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2012 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2013 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2014 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2015 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2016 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2017 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2018 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2019 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2020 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2021 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2022 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2023 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2024 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2025 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2026 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2027 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2028 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2029 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2030 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2031 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2032 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2033 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2034 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2035 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2036 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2037 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2038 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2039 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2040 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2041 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2042 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2043 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2044 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2045 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2046 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2047 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2048 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2049 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2050 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2051 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2052 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2053 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2054 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2055 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2056 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2057 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2058 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2059 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2060 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2061 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2062 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2063 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2064 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2065 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2066 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2067 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2068 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2069 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2070 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2071 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2072 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2073 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2074 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2075 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2076 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2077 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2078 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2079 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2080 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2081 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2082 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2083 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2084 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2085 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2086 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2087 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2088 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2089 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2090 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2091 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2092 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2093 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2094 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2095 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2096 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2097 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2098 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2099 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2100 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2101 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2102 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2103 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2104 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2105 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2106 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2107 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2108 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2109 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2110 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2111 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2112 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2113 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2114 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2115 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2116 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2117 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2118 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2119 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2120 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2121 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2122 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2123 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2124 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2125 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2126 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2127 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2128 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2129 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2130 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2131 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2132 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2133 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2134 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2135 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2136 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2137 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2138 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2139 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2140 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2141 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2142 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2143 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2144 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2145 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2146 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2147 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2148 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2149 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2150 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2151 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2152 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2153 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2154 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2155 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2156 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2157 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2158 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2159 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2160 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2161 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2162 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2163 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2164 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2165 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2166 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2167 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2168 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2169 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2170 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2171 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2172 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2173 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2174 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2175 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2176 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2177 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2178 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2179 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2180 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2181 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2182 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2183 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2184 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2185 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2186 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2187 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2188 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2189 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2190 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2191 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2192 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2193 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2194 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2195 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2196 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2197 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2198 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2199 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2200 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2201 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2202 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2203 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2204 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2205 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2206 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2207 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2208 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2209 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2210 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2211 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2212 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2213 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2214 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2215 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2216 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2217 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2218 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2219 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2220 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2221 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2222 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2223 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2224 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2225 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2226 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2227 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2228 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2229 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2230 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2231 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2232 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2233 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2234 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2235 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2236 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2237 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2238 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2239 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2240 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2241 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2242 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2243 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2244 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2245 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2246 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2247 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2248 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2249 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2250 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2251 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2252 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2253 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2254 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2255 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2256 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2257 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2258 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2259 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2260 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2261 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2262 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2263 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2264 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2265 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2266 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2267 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2268 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2269 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2270 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2271 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2272 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2273 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2274 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2275 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2276 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2277 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2278 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2279 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2280 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2281 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2282 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2283 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2284 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2285 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2286 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2287 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2288 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2289 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2290 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2291 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2292 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2293 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2294 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2295 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2296 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2297 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2298 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2299 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2300 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2301 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2302 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2303 VP V_da2_N outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2304 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2305 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2306 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2307 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2308 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2309 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2310 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2311 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2312 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2313 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2314 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2315 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2316 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2317 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2318 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2319 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2320 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2321 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2322 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2323 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2324 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2325 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2326 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2327 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2328 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2329 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2330 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2331 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2332 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2333 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2334 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2335 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2336 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2337 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2338 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2339 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2340 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2341 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2342 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2343 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2344 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2345 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2346 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2347 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2348 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2349 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2350 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2351 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2352 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2353 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2354 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2355 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2356 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2357 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2358 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2359 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2360 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2361 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2362 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2363 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2364 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2365 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2366 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2367 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2368 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2369 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2370 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2371 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2372 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2373 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2374 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2375 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2376 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2377 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2378 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2379 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2380 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2381 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2382 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2383 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2384 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2385 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2386 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2387 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2388 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2389 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2390 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2391 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2392 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2393 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2394 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2395 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2396 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2397 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2398 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2399 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2400 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2401 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2402 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2403 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2404 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2405 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2406 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2407 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2408 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2409 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2410 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2411 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2412 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2413 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2414 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2415 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2416 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2417 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2418 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2419 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2420 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2421 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2422 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2423 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2424 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2425 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2426 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2427 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2428 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2429 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2430 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2431 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2432 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2433 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2434 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2435 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2436 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2437 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2438 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2439 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2440 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2441 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2442 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2443 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2444 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2445 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2446 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2447 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2448 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2449 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2450 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2451 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2452 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2453 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2454 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2455 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2456 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2457 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2458 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2459 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2460 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2461 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2462 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2463 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2464 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2465 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2466 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2467 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2468 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2469 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2470 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2471 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2472 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2473 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2474 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2475 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2476 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2477 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2478 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2479 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2480 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2481 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2482 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2483 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2484 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2485 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2486 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2487 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2488 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2489 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2490 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2491 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2492 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2493 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2494 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2495 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2496 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2497 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2498 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2499 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2500 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2501 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2502 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2503 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2504 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2505 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2506 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2507 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2508 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2509 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2510 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2511 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2512 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2513 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2514 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2515 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2516 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2517 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2518 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2519 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2520 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2521 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2522 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2523 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2524 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2525 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2526 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2527 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2528 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2529 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2530 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2531 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2532 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2533 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2534 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2535 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2536 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2537 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2538 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2539 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2540 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2541 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2542 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2543 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2544 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2545 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2546 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2547 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2548 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2549 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2550 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2551 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2552 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2553 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2554 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2555 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2556 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2557 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2558 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2559 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2560 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2561 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2562 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2563 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2564 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2565 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2566 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2567 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2568 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2569 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2570 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2571 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2572 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2573 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2574 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2575 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2576 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2577 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2578 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2579 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2580 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2581 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2582 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2583 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2584 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2585 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2586 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2587 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2588 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2589 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2590 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2591 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2592 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2593 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2594 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2595 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2596 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2597 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2598 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2599 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2600 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2601 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2602 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2603 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2604 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2605 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2606 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2607 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2608 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2609 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2610 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2611 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2612 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2613 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2614 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2615 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2616 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2617 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2618 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2619 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2620 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2621 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2622 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2623 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2624 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2625 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2626 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2627 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2628 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2629 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2630 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2631 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2632 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2633 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2634 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2635 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2636 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2637 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2638 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2639 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2640 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2641 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2642 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2643 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2644 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2645 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2646 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2647 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2648 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2649 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2650 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2651 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2652 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2653 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2654 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2655 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2656 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2657 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2658 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2659 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2660 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2661 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2662 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2663 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2664 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2665 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2666 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2667 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2668 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2669 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2670 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2671 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2672 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2673 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2674 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2675 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2676 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2677 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2678 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2679 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2680 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2681 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2682 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2683 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2684 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2685 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2686 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2687 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2688 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2689 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2690 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2691 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2692 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2693 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2694 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2695 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2696 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2697 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2698 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2699 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2700 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2701 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2702 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2703 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2704 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2705 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2706 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2707 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2708 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2709 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2710 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2711 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2712 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2713 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2714 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2715 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2716 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2717 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2718 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2719 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2720 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2721 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2722 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2723 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2724 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2725 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2726 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2727 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2728 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2729 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2730 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2731 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2732 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2733 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2734 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2735 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2736 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2737 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2738 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2739 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2740 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2741 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2742 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2743 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2744 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2745 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2746 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2747 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2748 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2749 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2750 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2751 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2752 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2753 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2754 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2755 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2756 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2757 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2758 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2759 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2760 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2761 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2762 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2763 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2764 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2765 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2766 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2767 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2768 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2769 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2770 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2771 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2772 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2773 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2774 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2775 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2776 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2777 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2778 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2779 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2780 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2781 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2782 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2783 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2784 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2785 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2786 InputRef outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2787 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2788 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2789 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2790 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2791 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2792 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2793 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2794 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2795 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2796 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2797 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2798 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2799 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2800 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2801 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2802 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2803 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2804 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2805 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2806 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2807 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2808 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2809 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2810 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2811 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2812 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2813 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2814 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2815 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2816 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2817 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2818 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2819 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2820 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2821 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2822 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2823 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2824 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2825 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2826 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2827 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2828 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2829 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2830 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2831 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2832 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2833 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2834 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2835 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2836 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2837 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2838 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2839 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2840 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2841 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2842 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2843 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2844 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2845 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2846 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2847 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2848 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2849 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2850 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2851 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2852 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2853 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2854 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2855 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2856 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2857 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2858 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2859 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2860 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2861 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2862 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2863 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2864 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2865 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2866 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2867 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2868 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2869 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2870 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2871 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2872 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2873 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2874 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2875 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2876 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2877 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2878 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2879 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2880 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2881 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2882 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2883 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2884 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2885 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2886 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2887 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2888 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2889 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2890 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2891 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2892 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2893 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2894 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2895 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2896 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2897 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2898 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2899 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2900 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2901 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2902 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2903 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2904 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2905 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2906 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2907 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2908 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2909 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2910 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2911 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2912 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2913 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2914 V_da2_P VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2915 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2916 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2917 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2918 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2919 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2920 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2921 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2922 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2923 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2924 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2925 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2926 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2927 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2928 a_n19882_7120# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2929 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2930 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2931 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2932 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2933 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2934 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2935 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2936 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2937 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2938 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2939 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2940 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2941 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2942 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2943 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2944 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2945 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2946 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2947 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2948 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2949 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2950 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2951 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2952 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2953 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2954 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2955 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2956 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2957 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2958 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2959 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2960 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2961 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2962 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2963 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2964 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2965 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2966 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2967 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2968 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2969 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2970 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2971 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2972 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2973 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2974 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2975 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2976 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2977 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2978 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2979 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2980 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2981 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2982 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2983 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2984 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2985 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2986 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2987 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2988 VP V_da2_N outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X2989 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2990 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2991 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2992 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2993 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2994 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2995 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2996 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2997 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2998 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2999 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3000 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3001 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3002 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3003 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3004 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3005 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3006 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3007 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3008 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3009 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3010 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3011 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3012 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3013 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3014 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3015 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3016 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3017 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3018 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3019 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3020 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3021 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3022 V_da1_N VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3023 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3024 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3025 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3026 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3027 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3028 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3029 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3030 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3031 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3032 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3033 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3034 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3035 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3036 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3037 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3038 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3039 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3040 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3041 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3042 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3043 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3044 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3045 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3046 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3047 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3048 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3049 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3050 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3051 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3052 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3053 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3054 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3055 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3056 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3057 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3058 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3059 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3060 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3061 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3062 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3063 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3064 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3065 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3066 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3067 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3068 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3069 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3070 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3071 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3072 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3073 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3074 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3075 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3076 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3077 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3078 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3079 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3080 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3081 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3082 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3083 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3084 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3085 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3086 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3087 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3088 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3089 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3090 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3091 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3092 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3093 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3094 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3095 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3096 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3097 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3098 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3099 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3100 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3101 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3102 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3103 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3104 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3105 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3106 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3107 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3108 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3109 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3110 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3111 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3112 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3113 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3114 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3115 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3116 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3117 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3118 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3119 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3120 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3121 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3122 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3123 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3124 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3125 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3126 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3127 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3128 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3129 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3130 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3131 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3132 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3133 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3134 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3135 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3136 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3137 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3138 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3139 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3140 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3141 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3142 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3143 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3144 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3145 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3146 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3147 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3148 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3149 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3150 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3151 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3152 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3153 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3154 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3155 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3156 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3157 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3158 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3159 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3160 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3161 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3162 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3163 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3164 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3165 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3166 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3167 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3168 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3169 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3170 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3171 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3172 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3173 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3174 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3175 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3176 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3177 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3178 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3179 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3180 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3181 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3182 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3183 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3184 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3185 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3186 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3187 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3188 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3189 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3190 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3191 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3192 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3193 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3194 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3195 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3196 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3197 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3198 V_da1_P VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3199 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3200 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3201 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3202 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3203 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3204 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3205 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3206 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3207 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3208 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3209 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3210 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3211 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3212 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3213 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3214 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3215 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3216 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3217 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3218 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3219 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3220 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3221 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3222 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3223 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3224 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3225 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3226 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3227 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3228 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3229 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3230 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3231 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3232 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3233 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3234 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3235 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3236 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3237 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3238 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3239 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3240 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3241 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3242 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3243 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3244 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3245 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3246 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3247 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3248 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3249 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3250 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3251 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3252 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3253 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3254 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3255 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3256 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3257 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3258 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3259 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3260 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3261 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3262 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3263 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3264 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3265 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3266 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3267 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3268 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3269 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3270 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3271 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3272 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3273 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3274 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3275 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3276 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3277 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3278 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3279 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3280 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3281 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3282 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3283 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3284 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3285 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3286 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3287 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3288 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3289 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3290 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3291 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3292 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3293 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3294 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3295 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3296 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3297 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3298 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3299 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3300 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3301 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3302 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3303 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3304 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3305 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3306 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3307 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3308 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3309 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3310 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3311 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3312 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3313 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3314 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3315 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3316 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3317 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3318 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3319 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3320 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3321 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3322 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3323 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3324 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3325 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3326 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3327 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3328 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3329 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3330 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3331 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3332 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3333 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3334 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3335 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3336 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3337 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3338 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3339 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3340 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3341 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3342 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3343 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3344 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3345 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3346 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3347 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3348 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3349 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3350 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3351 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3352 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3353 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3354 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3355 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3356 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3357 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3358 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3359 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3360 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3361 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3362 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3363 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3364 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3365 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3366 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3367 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3368 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3369 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3370 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3371 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3372 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3373 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3374 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3375 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3376 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3377 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3378 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3379 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3380 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3381 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3382 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3383 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3384 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3385 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3386 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3387 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3388 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3389 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3390 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3391 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3392 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3393 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3394 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3395 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3396 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3397 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3398 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3399 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3400 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3401 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3402 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3403 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3404 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3405 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3406 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3407 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3408 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3409 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3410 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3411 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3412 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3413 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3414 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3415 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3416 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3417 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3418 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3419 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3420 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3421 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3422 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3423 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3424 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3425 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3426 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3427 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3428 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3429 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3430 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3431 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3432 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3433 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3434 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3435 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3436 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3437 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3438 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3439 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3440 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3441 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3442 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3443 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3444 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3445 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3446 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3447 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3448 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3449 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3450 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3451 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3452 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3453 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3454 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3455 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3456 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3457 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3458 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3459 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3460 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3461 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3462 InputRef outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3463 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3464 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3465 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3466 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3467 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3468 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3469 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3470 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3471 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3472 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3473 VP V_da2_P outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3474 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3475 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3476 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3477 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3478 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3479 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3480 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3481 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3482 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3483 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3484 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3485 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3486 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3487 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3488 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3489 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3490 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3491 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3492 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3493 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3494 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3495 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3496 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3497 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3498 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3499 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3500 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3501 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3502 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3503 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3504 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3505 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3506 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3507 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3508 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3509 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3510 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3511 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3512 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3513 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3514 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3515 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3516 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3517 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3518 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3519 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3520 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3521 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3522 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3523 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3524 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3525 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3526 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3527 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3528 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3529 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3530 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3531 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3532 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3533 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3534 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3535 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3536 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3537 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3538 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3539 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3540 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3541 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3542 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3543 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3544 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3545 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3546 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3547 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3548 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3549 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3550 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3551 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3552 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3553 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3554 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3555 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3556 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3557 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3558 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3559 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3560 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3561 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3562 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3563 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3564 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3565 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3566 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3567 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3568 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3569 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3570 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3571 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3572 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3573 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3574 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3575 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3576 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3577 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3578 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3579 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3580 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3581 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3582 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3583 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3584 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3585 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3586 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3587 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3588 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3589 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3590 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3591 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3592 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3593 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3594 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3595 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3596 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3597 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3598 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3599 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3600 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3601 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3602 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3603 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3604 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3605 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3606 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3607 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3608 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3609 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3610 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3611 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3612 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3613 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3614 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3615 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3616 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3617 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3618 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3619 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3620 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3621 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3622 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3623 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3624 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3625 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3626 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3627 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3628 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3629 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3630 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3631 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3632 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3633 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3634 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3635 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3636 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3637 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3638 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3639 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3640 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3641 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3642 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3643 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3644 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3645 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3646 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3647 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3648 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3649 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3650 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3651 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3652 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3653 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3654 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3655 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3656 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3657 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3658 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3659 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3660 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3661 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3662 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3663 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3664 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3665 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3666 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3667 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3668 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3669 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3670 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3671 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3672 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3673 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3674 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3675 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3676 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3677 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3678 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3679 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3680 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3681 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3682 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3683 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3684 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3685 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3686 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3687 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3688 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3689 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3690 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3691 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3692 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3693 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3694 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3695 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3696 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3697 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3698 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3699 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3700 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3701 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3702 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3703 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3704 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3705 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3706 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3707 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3708 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3709 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3710 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3711 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3712 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3713 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3714 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3715 V_da1_P VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3716 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3717 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3718 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3719 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3720 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3721 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3722 V_da1_N VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3723 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3724 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3725 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3726 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3727 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3728 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3729 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3730 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3731 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3732 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3733 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3734 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3735 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3736 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3737 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3738 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3739 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3740 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3741 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3742 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3743 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3744 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3745 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3746 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3747 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3748 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3749 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3750 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3751 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3752 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3753 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3754 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3755 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3756 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3757 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3758 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3759 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3760 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3761 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3762 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3763 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3764 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3765 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3766 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3767 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3768 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3769 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3770 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3771 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3772 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3773 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3774 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3775 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3776 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3777 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3778 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3779 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3780 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3781 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3782 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3783 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3784 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3785 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3786 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3787 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3788 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3789 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3790 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3791 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3792 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3793 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3794 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3795 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3796 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3797 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3798 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3799 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3800 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3801 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3802 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3803 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3804 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3805 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3806 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3807 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3808 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3809 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3810 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3811 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3812 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3813 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3814 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3815 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3816 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3817 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3818 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3819 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3820 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3821 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3822 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3823 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3824 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3825 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3826 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3827 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3828 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3829 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3830 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3831 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3832 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3833 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3834 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3835 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3836 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3837 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3838 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3839 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3840 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3841 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3842 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3843 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3844 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3845 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3846 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3847 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3848 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3849 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3850 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3851 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3852 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3853 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3854 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3855 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3856 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3857 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3858 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3859 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3860 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3861 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3862 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3863 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3864 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3865 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3866 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3867 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3868 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3869 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3870 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3871 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3872 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3873 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3874 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3875 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3876 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3877 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3878 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3879 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3880 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3881 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3882 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3883 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3884 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3885 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3886 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3887 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3888 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3889 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3890 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3891 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3892 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3893 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3894 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3895 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3896 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3897 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3898 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3899 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3900 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3901 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3902 VP V_da2_P outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X3903 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3904 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3905 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3906 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3907 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3908 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3909 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3910 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3911 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3912 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3913 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3914 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3915 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3916 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3917 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3918 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3919 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3920 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3921 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3922 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3923 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3924 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3925 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3926 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3927 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3928 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3929 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3930 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3931 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3932 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3933 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3934 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3935 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3936 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3937 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3938 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3939 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3940 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3941 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3942 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3943 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3944 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3945 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3946 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3947 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3948 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3949 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3950 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3951 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3952 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3953 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3954 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3955 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3956 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3957 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3958 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3959 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3960 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3961 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3962 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3963 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3964 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3965 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3966 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3967 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3968 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3969 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3970 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19882_7120# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3971 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3972 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3973 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3974 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3975 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3976 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3977 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3978 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3979 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3980 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3981 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3982 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3983 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3984 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3985 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3986 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3987 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3988 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3989 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3990 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3991 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3992 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3993 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3994 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3995 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3996 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3997 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3998 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3999 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4000 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4001 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4002 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4003 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4004 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4005 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4006 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4007 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4008 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4009 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4010 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4011 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4012 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4013 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4014 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4015 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4016 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4017 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4018 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4019 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4020 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4021 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4022 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4023 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4024 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4025 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4026 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4027 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4028 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4029 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4030 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4031 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4032 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4033 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4034 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4035 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4036 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4037 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4038 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4039 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4040 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4041 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4042 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4043 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4044 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4045 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4046 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4047 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4048 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4049 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4050 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4051 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4052 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4053 V_da2_N VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4054 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4055 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4056 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4057 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4058 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4059 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4060 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4061 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4062 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4063 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4064 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4065 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4066 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4067 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4068 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4069 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4070 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4071 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4072 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4073 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4074 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4075 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4076 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4077 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4078 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4079 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4080 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4081 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4082 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4083 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4084 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4085 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4086 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4087 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4088 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4089 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4090 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4091 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4092 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4093 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4094 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4095 VP V_da2_N outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4096 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4097 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4098 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4099 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4100 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4101 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4102 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4103 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4104 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4105 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4106 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4107 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4108 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4109 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4110 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4111 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4112 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4113 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4114 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4115 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4116 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4117 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4118 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4119 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4120 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4121 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4122 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4123 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4124 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4125 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4126 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4127 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4128 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4129 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4130 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4131 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4132 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4133 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4134 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4135 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4136 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4137 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4138 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4139 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4140 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4141 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4142 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4143 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4144 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4145 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4146 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4147 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4148 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4149 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4150 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4151 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4152 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4153 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4154 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4155 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4156 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4157 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4158 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4159 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4160 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4161 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4162 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4163 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4164 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4165 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4166 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4167 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4168 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4169 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4170 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4171 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4172 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4173 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4174 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4175 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4176 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4177 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4178 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4179 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4180 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4181 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4182 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4183 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4184 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4185 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4186 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4187 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4188 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4189 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4190 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4191 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4192 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4193 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4194 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4195 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4196 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4197 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4198 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4199 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4200 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4201 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4202 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4203 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4204 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4205 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4206 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4207 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4208 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4209 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4210 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4211 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4212 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4213 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4214 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4215 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4216 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4217 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4218 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4219 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4220 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4221 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4222 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4223 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4224 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4225 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4226 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4227 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4228 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4229 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4230 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4231 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4232 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4233 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4234 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4235 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4236 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4237 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4238 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4239 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4240 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4241 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4242 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4243 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4244 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4245 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4246 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4247 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4248 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4249 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4250 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4251 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4252 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4253 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4254 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4255 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4256 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4257 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4258 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4259 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4260 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4261 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4262 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4263 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4264 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4265 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4266 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4267 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4268 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4269 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4270 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4271 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4272 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4273 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4274 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4275 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4276 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4277 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4278 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4279 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4280 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4281 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4282 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4283 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4284 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4285 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4286 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4287 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4288 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4289 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4290 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4291 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4292 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4293 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4294 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4295 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4296 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4297 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4298 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4299 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4300 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4301 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4302 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4303 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4304 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4305 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4306 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4307 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4308 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4309 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4310 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4311 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4312 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4313 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4314 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4315 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4316 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4317 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4318 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4319 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4320 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4321 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4322 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4323 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4324 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4325 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4326 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4327 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4328 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4329 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4330 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4331 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4332 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4333 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4334 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4335 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4336 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4337 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4338 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4339 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4340 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4341 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4342 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4343 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4344 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4345 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4346 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4347 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4348 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4349 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4350 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4351 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4352 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4353 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4354 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4355 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4356 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4357 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4358 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4359 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4360 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4361 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4362 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4363 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4364 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4365 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4366 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4367 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4368 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4369 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4370 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4371 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4372 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4373 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4374 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4375 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4376 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4377 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4378 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4379 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4380 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4381 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4382 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4383 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4384 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4385 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4386 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4387 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4388 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4389 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4390 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4391 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4392 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4393 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4394 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4395 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4396 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4397 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4398 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4399 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4400 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4401 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4402 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4403 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4404 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4405 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4406 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4407 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4408 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4409 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4410 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4411 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4412 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4413 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4414 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4415 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4416 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4417 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4418 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4419 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4420 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4421 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4422 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4423 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4424 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4425 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4426 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4427 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4428 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4429 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4430 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4431 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4432 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4433 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4434 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4435 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4436 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4437 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4438 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4439 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4440 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4441 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4442 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4443 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4444 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4445 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4446 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4447 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4448 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4449 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4450 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4451 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4452 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4453 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4454 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4455 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4456 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4457 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4458 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4459 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4460 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4461 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4462 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4463 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4464 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4465 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4466 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4467 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4468 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4469 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4470 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4471 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4472 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4473 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4474 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4475 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4476 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4477 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4478 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4479 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4480 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4481 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4482 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4483 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4484 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4485 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4486 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4487 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4488 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4489 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4490 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4491 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4492 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4493 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4494 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4495 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4496 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4497 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4498 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4499 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4500 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4501 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4502 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4503 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4504 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4505 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4506 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4507 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4508 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4509 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4510 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4511 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4512 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4513 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4514 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4515 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4516 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4517 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4518 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4519 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4520 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4521 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4522 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4523 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4524 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4525 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4526 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4527 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4528 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4529 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4530 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4531 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4532 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4533 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4534 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4535 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4536 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4537 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4538 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4539 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4540 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4541 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4542 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4543 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4544 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4545 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4546 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4547 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4548 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4549 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4550 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4551 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4552 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4553 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4554 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4555 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4556 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4557 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4558 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4559 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4560 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4561 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4562 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4563 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4564 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4565 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4566 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4567 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4568 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4569 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4570 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4571 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4572 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4573 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4574 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4575 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4576 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4577 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4578 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4579 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4580 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4581 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4582 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4583 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4584 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4585 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4586 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4587 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4588 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4589 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4590 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4591 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4592 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4593 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4594 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4595 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4596 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4597 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4598 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4599 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4600 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4601 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4602 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4603 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4604 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4605 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4606 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4607 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4608 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4609 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4610 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4611 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4612 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4613 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4614 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4615 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4616 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4617 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4618 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4619 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4620 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4621 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4622 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4623 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4624 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4625 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4626 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4627 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4628 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4629 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4630 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4631 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4632 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4633 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4634 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4635 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4636 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4637 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4638 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4639 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4640 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4641 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4642 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4643 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4644 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4645 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4646 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4647 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4648 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4649 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4650 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4651 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4652 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4653 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4654 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4655 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4656 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4657 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4658 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4659 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4660 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4661 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4662 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4663 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4664 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4665 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4666 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4667 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4668 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4669 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4670 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4671 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4672 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4673 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4674 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4675 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4676 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4677 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4678 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4679 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4680 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4681 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4682 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4683 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4684 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4685 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4686 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4687 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4688 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4689 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4690 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4691 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4692 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4693 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4694 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4695 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4696 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4697 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4698 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4699 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4700 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4701 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4702 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4703 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4704 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4705 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4706 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4707 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4708 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4709 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4710 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4711 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4712 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4713 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4714 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4715 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4716 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4717 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4718 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4719 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4720 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4721 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4722 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4723 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4724 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4725 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4726 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4727 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4728 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4729 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4730 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4731 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4732 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4733 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4734 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4735 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4736 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4737 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4738 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4739 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4740 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4741 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4742 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4743 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4744 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4745 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4746 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4747 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4748 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4749 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4750 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4751 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4752 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4753 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4754 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4755 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4756 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4757 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4758 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4759 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4760 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4761 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4762 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4763 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4764 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4765 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4766 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4767 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4768 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4769 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4770 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4771 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4772 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4773 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4774 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4775 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4776 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4777 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4778 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4779 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4780 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4781 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4782 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4783 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4784 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4785 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4786 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4787 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4788 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4789 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4790 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4791 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4792 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4793 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4794 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4795 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4796 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4797 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4798 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4799 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4800 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4801 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4802 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4803 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4804 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4805 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4806 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4807 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4808 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4809 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4810 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4811 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4812 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4813 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4814 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4815 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4816 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4817 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4818 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4819 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4820 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4821 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4822 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4823 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4824 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4825 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4826 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4827 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4828 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4829 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4830 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4831 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4832 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4833 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4834 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4835 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4836 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4837 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4838 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4839 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4840 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4841 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4842 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4843 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4844 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4845 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4846 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4847 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4848 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4849 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4850 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4851 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4852 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4853 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4854 I_Bias I_Bias a_n19882_7120# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4855 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4856 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4857 outd_stage3_0/outd_stage2_0/VN I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X4858 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4859 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4860 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4861 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4862 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4863 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4864 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4865 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4866 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4867 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4868 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4869 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4870 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4871 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4872 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4873 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4874 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4875 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4876 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4877 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4878 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4879 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4880 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4881 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4882 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4883 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4884 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4885 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4886 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4887 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4888 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4889 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4890 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4891 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4892 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4893 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4894 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4895 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4896 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4897 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4898 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4899 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4900 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4901 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4902 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4903 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4904 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4905 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4906 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4907 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4908 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4909 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4910 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4911 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4912 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4913 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4914 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4915 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4916 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4917 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4918 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4919 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4920 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4921 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4922 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4923 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4924 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4925 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4926 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4927 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4928 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4929 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4930 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4931 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4932 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4933 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4934 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4935 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4936 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4937 outd_stage3_0/outd_stage2_0/VN I_Bias sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X4938 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4939 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4940 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4941 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X4942 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4943 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4944 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4945 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4946 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4947 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4948 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4949 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4950 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4951 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4952 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4953 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4954 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4955 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4956 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4957 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4958 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4959 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4960 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4961 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4962 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4963 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4964 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4965 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4966 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4967 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4968 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4969 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4970 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4971 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4972 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4973 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4974 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4975 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4976 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4977 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4978 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4979 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4980 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4981 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4982 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4983 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4984 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4985 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4986 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4987 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4988 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4989 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4990 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4991 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4992 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4993 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4994 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4995 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4996 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4997 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4998 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4999 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5000 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5001 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5002 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5003 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5004 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5005 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5006 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5007 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5008 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5009 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5010 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5011 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5012 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5013 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5014 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5015 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5016 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5017 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5018 V_da2_P VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5019 outd_stage1_0/isource_out InputRef V_da1_N outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5020 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5021 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5022 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5023 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5024 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5025 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5026 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5027 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5028 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5029 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5030 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5031 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5032 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5033 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5034 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5035 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5036 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5037 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5038 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5039 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5040 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5041 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5042 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5043 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5044 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5045 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5046 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5047 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5048 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5049 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5050 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5051 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5052 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5053 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5054 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5055 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5056 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5057 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5058 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5059 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5060 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5061 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5062 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5063 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5064 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5065 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5066 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5067 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5068 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5069 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5070 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5071 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5072 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5073 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5074 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5075 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5076 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5077 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5078 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5079 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5080 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5081 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5082 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5083 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5084 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5085 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5086 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5087 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5088 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5089 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5090 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5091 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5092 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5093 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5094 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5095 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5096 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5097 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5098 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5099 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5100 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5101 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5102 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5103 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5104 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5105 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5106 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5107 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5108 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5109 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5110 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5111 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5112 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5113 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5114 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5115 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5116 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5117 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5118 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5119 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5120 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5121 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5122 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5123 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5124 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5125 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5126 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5127 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5128 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5129 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5130 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5131 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5132 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5133 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5134 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5135 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5136 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5137 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5138 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5139 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5140 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5141 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5142 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5143 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5144 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5145 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5146 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5147 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5148 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5149 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5150 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5151 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5152 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5153 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5154 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5155 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5156 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5157 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5158 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5159 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5160 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5161 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5162 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5163 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5164 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5165 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5166 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5167 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5168 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5169 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5170 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5171 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5172 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5173 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5174 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5175 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5176 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5177 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5178 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5179 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5180 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5181 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5182 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5183 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5184 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5185 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5186 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5187 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5188 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5189 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5190 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5191 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5192 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5193 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5194 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5195 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5196 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5197 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5198 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5199 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5200 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5201 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5202 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5203 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5204 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5205 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5206 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5207 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5208 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5209 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5210 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5211 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5212 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5213 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5214 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5215 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5216 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5217 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5218 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5219 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5220 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5221 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5222 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5223 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5224 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5225 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5226 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5227 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5228 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5229 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5230 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5231 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5232 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5233 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5234 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5235 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5236 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5237 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5238 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5239 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5240 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5241 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5242 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5243 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5244 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5245 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5246 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5247 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5248 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5249 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5250 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5251 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5252 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5253 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5254 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5255 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5256 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5257 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5258 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5259 outd_stage3_0/outd_stage2_0/VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5260 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5261 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5262 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5263 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5264 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5265 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5266 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5267 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5268 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5269 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5270 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5271 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5272 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5273 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5274 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5275 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5276 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5277 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5278 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5279 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5280 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5281 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5282 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5283 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5284 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5285 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5286 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5287 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5288 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5289 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5290 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5291 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5292 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5293 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5294 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5295 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5296 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5297 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5298 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5299 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5300 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5301 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5302 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5303 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5304 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5305 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5306 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5307 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5308 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5309 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5310 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5311 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5312 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5313 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5314 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5315 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5316 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5317 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5318 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5319 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5320 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5321 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5322 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5323 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5324 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5325 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5326 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5327 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5328 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5329 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5330 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5331 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5332 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5333 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5334 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5335 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5336 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5337 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5338 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5339 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5340 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5341 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5342 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5343 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5344 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5345 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5346 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5347 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5348 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5349 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5350 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5351 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5352 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5353 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5354 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5355 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5356 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5357 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5358 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5359 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5360 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5361 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5362 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5363 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5364 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5365 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5366 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5367 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5368 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5369 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5370 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5371 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5372 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5373 a_n19882_7120# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5374 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5375 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5376 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5377 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5378 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5379 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5380 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5381 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5382 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5383 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5384 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5385 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5386 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5387 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5388 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5389 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5390 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5391 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5392 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5393 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5394 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5395 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5396 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5397 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5398 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5399 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5400 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5401 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5402 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5403 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5404 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5405 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5406 OutputN VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5407 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5408 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5409 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5410 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5411 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5412 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5413 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5414 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5415 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5416 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5417 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5418 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5419 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5420 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5421 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5422 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5423 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5424 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5425 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5426 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5427 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5428 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5429 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5430 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5431 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5432 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5433 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5434 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5435 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5436 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5437 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5438 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5439 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5440 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5441 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5442 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5443 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5444 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5445 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5446 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5447 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5448 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5449 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5450 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5451 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5452 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5453 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5454 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5455 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5456 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5457 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5458 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5459 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5460 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5461 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5462 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5463 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5464 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5465 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5466 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5467 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5468 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5469 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5470 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5471 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5472 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5473 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5474 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5475 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5476 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5477 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5478 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5479 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5480 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5481 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5482 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5483 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5484 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5485 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5486 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5487 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5488 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5489 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5490 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5491 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5492 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5493 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5494 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5495 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5496 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5497 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5498 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5499 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5500 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5501 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5502 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5503 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5504 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5505 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5506 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5507 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5508 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5509 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5510 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5511 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5512 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5513 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5514 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5515 V_da1_N InputRef outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5516 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5517 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5518 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5519 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5520 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5521 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5522 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5523 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5524 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5525 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5526 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5527 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5528 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5529 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5530 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5531 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5532 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5533 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5534 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5535 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5536 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5537 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5538 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5539 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5540 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5541 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5542 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5543 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5544 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5545 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5546 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5547 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5548 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5549 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5550 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5551 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5552 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5553 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5554 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5555 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5556 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5557 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5558 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5559 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5560 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5561 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5562 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5563 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5564 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5565 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5566 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5567 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5568 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5569 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5570 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5571 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5572 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5573 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5574 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5575 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5576 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5577 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5578 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5579 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5580 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5581 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5582 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5583 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5584 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5585 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5586 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5587 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5588 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5589 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5590 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5591 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5592 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5593 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5594 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5595 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5596 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5597 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5598 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5599 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5600 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5601 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5602 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5603 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5604 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5605 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5606 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5607 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5608 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5609 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5610 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5611 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5612 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5613 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5614 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5615 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5616 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5617 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5618 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5619 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5620 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5621 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5622 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5623 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5624 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5625 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5626 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5627 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5628 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5629 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5630 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5631 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5632 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5633 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5634 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5635 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5636 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5637 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5638 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5639 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5640 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5641 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5642 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5643 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5644 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5645 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5646 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5647 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5648 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5649 V_da2_N VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5650 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5651 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5652 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5653 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5654 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5655 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5656 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5657 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5658 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5659 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5660 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5661 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5662 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5663 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5664 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5665 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5666 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5667 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5668 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5669 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5670 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5671 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5672 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5673 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5674 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5675 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5676 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5677 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5678 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5679 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5680 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5681 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5682 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5683 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5684 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5685 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5686 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5687 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5688 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5689 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5690 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5691 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5692 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5693 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5694 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5695 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5696 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5697 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5698 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5699 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5700 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5701 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5702 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5703 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5704 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5705 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5706 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5707 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5708 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5709 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5710 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5711 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5712 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5713 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5714 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5715 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5716 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5717 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5718 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5719 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5720 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5721 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5722 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5723 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5724 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5725 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5726 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5727 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5728 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5729 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5730 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5731 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5732 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5733 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5734 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5735 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5736 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5737 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5738 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5739 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5740 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5741 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5742 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5743 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5744 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5745 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5746 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5747 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5748 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5749 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5750 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5751 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5752 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5753 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5754 VP V_da2_P outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5755 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5756 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5757 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5758 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5759 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5760 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5761 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5762 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5763 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5764 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5765 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5766 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5767 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5768 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5769 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5770 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5771 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5772 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5773 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5774 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5775 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5776 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5777 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5778 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5779 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5780 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5781 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5782 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5783 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5784 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5785 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5786 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5787 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5788 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5789 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5790 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5791 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5792 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5793 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5794 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5795 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5796 V_da2_N V_da1_N outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5797 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5798 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5799 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5800 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5801 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5802 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5803 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5804 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5805 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5806 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5807 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5808 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5809 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5810 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5811 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5812 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5813 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5814 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5815 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5816 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5817 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5818 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5819 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5820 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5821 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5822 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5823 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5824 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5825 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5826 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5827 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5828 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5829 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5830 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5831 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5832 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5833 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5834 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5835 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5836 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5837 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5838 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5839 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5840 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5841 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5842 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5843 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5844 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5845 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5846 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5847 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5848 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5849 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5850 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5851 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5852 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5853 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5854 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5855 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5856 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5857 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5858 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5859 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5860 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5861 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5862 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5863 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5864 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5865 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5866 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5867 VP OutputN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5868 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5869 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5870 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5871 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5872 a_n19260_7126# I_Bias outd_stage1_0/isource_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5873 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5874 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5875 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5876 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5877 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5878 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5879 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5880 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5881 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5882 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5883 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5884 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5885 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5886 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5887 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5888 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5889 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5890 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5891 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5892 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5893 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5894 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5895 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5896 V_da2_P V_da1_P outd_stage2_0/cmirror_out outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5897 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5898 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5899 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5900 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5901 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5902 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5903 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5904 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5905 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5906 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5907 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5908 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5909 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5910 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5911 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5912 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5913 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5914 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5915 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5916 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5917 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5918 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5919 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5920 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5921 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5922 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5923 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5924 V_da1_P InputSignal outd_stage1_0/isource_out outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5925 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5926 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5927 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5928 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5929 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5930 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5931 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5932 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5933 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5934 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5935 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5936 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5937 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5938 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5939 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5940 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5941 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5942 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5943 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5944 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5945 VP OutputP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X5946 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5947 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5948 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5949 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5950 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5951 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5952 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5953 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5954 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5955 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5956 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5957 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5958 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5959 OutputN V_da2_N outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5960 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5961 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5962 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5963 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5964 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5965 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5966 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5967 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5968 outd_stage1_0/isource_out InputSignal V_da1_P outd_stage1_0/isource_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5969 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5970 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5971 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5972 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5973 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5974 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5975 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5976 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5977 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5978 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_N OutputN outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5979 outd_stage3_0/outd_stage2_0/cmirror_out V_da2_P OutputP outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5980 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5981 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5982 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5983 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5984 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5985 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5986 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5987 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5988 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5989 OutputP V_da2_P outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5990 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5991 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5992 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5993 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5994 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5995 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X5996 outd_stage2_0/cmirror_out V_da1_P V_da2_P outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5997 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5998 a_n14090_6326# I_Bias outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5999 outd_stage3_0/outd_stage2_0/VN I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6000 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6001 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6002 OutputP VP outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__res_high_po_5p73 l=4e+06u
X6003 outd_stage1_0/isource_out I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6004 a_n14090_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6005 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6006 a_n19260_7126# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6007 outd_stage2_0/cmirror_out I_Bias a_n14090_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6008 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6009 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/cmirror_out outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6010 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6011 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6012 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6013 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6014 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6015 outd_stage2_0/cmirror_out V_da1_N V_da2_N outd_stage2_0/cmirror_out sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6016 outd_stage3_0/outd_stage2_0/VN I_Bias a_n19260_7126# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6017 a_230_6326# I_Bias outd_stage3_0/outd_stage2_0/VN outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6018 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6019 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X6020 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6021 outd_stage3_0/outd_stage2_0/cmirror_out I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6022 outd_stage3_0/outd_stage2_0/VN I_Bias a_230_6326# outd_stage3_0/outd_stage2_0/VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
