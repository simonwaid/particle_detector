magic
tech sky130B
magscale 1 2
timestamp 1654683408
<< pwell >>
rect 130 1200 1498 1266
rect 132 740 1498 756
rect 132 706 1500 740
rect 132 690 1498 706
rect 132 632 1498 648
rect 132 598 1500 632
rect 132 582 1498 598
rect 132 72 1498 138
<< poly >>
rect 130 1200 1498 1266
rect 132 740 1498 756
rect 132 706 1500 740
rect 132 690 1498 706
rect 132 632 1498 648
rect 132 598 1500 632
rect 132 582 1498 598
rect 132 72 1498 138
<< locali >>
rect 130 1216 1498 1250
rect 132 706 1500 740
rect 132 598 1500 632
rect 132 88 1498 122
<< metal1 >>
rect 70 1210 1560 1260
rect 188 1002 198 1178
rect 252 1002 262 1178
rect 424 1002 434 1178
rect 488 1002 498 1178
rect 660 1002 670 1178
rect 724 1002 734 1178
rect 896 1002 906 1178
rect 960 1002 970 1178
rect 1132 1002 1142 1178
rect 1196 1002 1206 1178
rect 1368 1002 1378 1178
rect 1432 1002 1442 1178
rect 70 778 80 954
rect 134 778 144 954
rect 306 778 316 954
rect 370 778 380 954
rect 542 778 552 954
rect 606 778 616 954
rect 778 778 788 954
rect 842 778 852 954
rect 1014 778 1024 954
rect 1078 778 1088 954
rect 1250 778 1260 954
rect 1314 778 1324 954
rect 1486 778 1496 954
rect 1550 778 1560 954
rect 70 700 1560 750
rect 70 590 1560 640
rect 188 384 198 560
rect 252 384 262 560
rect 424 384 434 560
rect 488 384 498 560
rect 660 384 670 560
rect 724 384 734 560
rect 896 384 906 560
rect 960 384 970 560
rect 1132 384 1142 560
rect 1196 384 1206 560
rect 1368 384 1378 560
rect 1432 384 1442 560
rect 70 160 80 336
rect 134 160 144 336
rect 306 160 316 336
rect 370 160 380 336
rect 542 160 552 336
rect 606 160 616 336
rect 778 160 788 336
rect 842 160 852 336
rect 1014 160 1024 336
rect 1078 160 1088 336
rect 1250 160 1260 336
rect 1314 160 1324 336
rect 1486 160 1496 336
rect 1550 160 1560 336
rect 70 80 1560 130
<< via1 >>
rect 198 1002 252 1178
rect 434 1002 488 1178
rect 670 1002 724 1178
rect 906 1002 960 1178
rect 1142 1002 1196 1178
rect 1378 1002 1432 1178
rect 80 778 134 954
rect 316 778 370 954
rect 552 778 606 954
rect 788 778 842 954
rect 1024 778 1078 954
rect 1260 778 1314 954
rect 1496 778 1550 954
rect 198 384 252 560
rect 434 384 488 560
rect 670 384 724 560
rect 906 384 960 560
rect 1142 384 1196 560
rect 1378 384 1432 560
rect 80 160 134 336
rect 316 160 370 336
rect 552 160 606 336
rect 788 160 842 336
rect 1024 160 1078 336
rect 1260 160 1314 336
rect 1496 160 1550 336
<< metal2 >>
rect 190 1178 1440 1190
rect 190 1030 198 1178
rect 252 1030 434 1178
rect 198 992 252 1002
rect 488 1030 670 1178
rect 434 992 488 1002
rect 724 1030 906 1178
rect 670 992 724 1002
rect 960 1030 1142 1178
rect 906 992 960 1002
rect 1196 1030 1378 1178
rect 1142 992 1196 1002
rect 1432 1030 1440 1178
rect 1378 992 1432 1002
rect 80 954 134 964
rect 70 778 80 920
rect 316 954 370 964
rect 134 778 316 920
rect 552 954 606 964
rect 370 778 552 920
rect 788 954 842 964
rect 606 778 788 920
rect 1024 954 1078 964
rect 842 778 1024 920
rect 1260 954 1314 964
rect 1078 778 1260 920
rect 1496 954 1550 964
rect 1314 778 1496 920
rect 1550 778 1560 920
rect 70 760 1560 778
rect 190 560 1440 570
rect 190 410 198 560
rect 252 410 434 560
rect 198 374 252 384
rect 488 410 670 560
rect 434 374 488 384
rect 724 410 906 560
rect 670 374 724 384
rect 960 410 1142 560
rect 906 374 960 384
rect 1196 410 1378 560
rect 1142 374 1196 384
rect 1432 410 1440 560
rect 1378 374 1432 384
rect 80 336 134 346
rect 70 160 80 300
rect 316 336 370 346
rect 134 160 316 300
rect 552 336 606 346
rect 370 160 552 300
rect 788 336 842 346
rect 606 160 788 300
rect 1024 336 1078 346
rect 842 160 1024 300
rect 1260 336 1314 346
rect 1078 160 1260 300
rect 1496 336 1550 346
rect 1314 160 1496 300
rect 1550 160 1560 300
rect 70 140 1560 160
use sky130_fd_pr__nfet_01v8_lvt_ZHX6G9  sky130_fd_pr__nfet_01v8_lvt_ZHX6G9_0
timestamp 1654683408
transform 1 0 815 0 1 669
box -875 -719 875 719
<< end >>
