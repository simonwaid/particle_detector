magic
tech sky130A
magscale 1 2
timestamp 1645802395
<< metal3 >>
rect -1350 1072 1349 1100
rect -1350 -1072 1265 1072
rect 1329 -1072 1349 1072
rect -1350 -1100 1349 -1072
<< via3 >>
rect 1265 -1072 1329 1072
<< mimcap >>
rect -1250 960 1150 1000
rect -1250 -960 -1210 960
rect 1110 -960 1150 960
rect -1250 -1000 1150 -960
<< mimcapcontact >>
rect -1210 -960 1110 960
<< metal4 >>
rect 1249 1072 1345 1088
rect -1211 960 1111 961
rect -1211 -960 -1210 960
rect 1110 -960 1111 960
rect -1211 -961 1111 -960
rect 1249 -1072 1265 1072
rect 1329 -1072 1345 1072
rect 1249 -1088 1345 -1072
<< properties >>
string FIXED_BBOX -1350 -1100 1250 1100
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 12 l 10 val 248.36 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
