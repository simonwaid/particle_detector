magic
tech sky130A
magscale 1 2
timestamp 1645781187
<< error_p >>
rect -617 272 -559 278
rect -421 272 -363 278
rect -225 272 -167 278
rect -29 272 29 278
rect 167 272 225 278
rect 363 272 421 278
rect 559 272 617 278
rect -617 238 -605 272
rect -421 238 -409 272
rect -225 238 -213 272
rect -29 238 -17 272
rect 167 238 179 272
rect 363 238 375 272
rect 559 238 571 272
rect -617 232 -559 238
rect -421 232 -363 238
rect -225 232 -167 238
rect -29 232 29 238
rect 167 232 225 238
rect 363 232 421 238
rect 559 232 617 238
rect -715 -238 -657 -232
rect -519 -238 -461 -232
rect -323 -238 -265 -232
rect -127 -238 -69 -232
rect 69 -238 127 -232
rect 265 -238 323 -232
rect 461 -238 519 -232
rect 657 -238 715 -232
rect -715 -272 -703 -238
rect -519 -272 -507 -238
rect -323 -272 -311 -238
rect -127 -272 -115 -238
rect 69 -272 81 -238
rect 265 -272 277 -238
rect 461 -272 473 -238
rect 657 -272 669 -238
rect -715 -278 -657 -272
rect -519 -278 -461 -272
rect -323 -278 -265 -272
rect -127 -278 -69 -272
rect 69 -278 127 -272
rect 265 -278 323 -272
rect 461 -278 519 -272
rect 657 -278 715 -272
<< pwell >>
rect -902 -410 902 410
<< nmos >>
rect -706 -200 -666 200
rect -608 -200 -568 200
rect -510 -200 -470 200
rect -412 -200 -372 200
rect -314 -200 -274 200
rect -216 -200 -176 200
rect -118 -200 -78 200
rect -20 -200 20 200
rect 78 -200 118 200
rect 176 -200 216 200
rect 274 -200 314 200
rect 372 -200 412 200
rect 470 -200 510 200
rect 568 -200 608 200
rect 666 -200 706 200
<< ndiff >>
rect -764 188 -706 200
rect -764 -188 -752 188
rect -718 -188 -706 188
rect -764 -200 -706 -188
rect -666 188 -608 200
rect -666 -188 -654 188
rect -620 -188 -608 188
rect -666 -200 -608 -188
rect -568 188 -510 200
rect -568 -188 -556 188
rect -522 -188 -510 188
rect -568 -200 -510 -188
rect -470 188 -412 200
rect -470 -188 -458 188
rect -424 -188 -412 188
rect -470 -200 -412 -188
rect -372 188 -314 200
rect -372 -188 -360 188
rect -326 -188 -314 188
rect -372 -200 -314 -188
rect -274 188 -216 200
rect -274 -188 -262 188
rect -228 -188 -216 188
rect -274 -200 -216 -188
rect -176 188 -118 200
rect -176 -188 -164 188
rect -130 -188 -118 188
rect -176 -200 -118 -188
rect -78 188 -20 200
rect -78 -188 -66 188
rect -32 -188 -20 188
rect -78 -200 -20 -188
rect 20 188 78 200
rect 20 -188 32 188
rect 66 -188 78 188
rect 20 -200 78 -188
rect 118 188 176 200
rect 118 -188 130 188
rect 164 -188 176 188
rect 118 -200 176 -188
rect 216 188 274 200
rect 216 -188 228 188
rect 262 -188 274 188
rect 216 -200 274 -188
rect 314 188 372 200
rect 314 -188 326 188
rect 360 -188 372 188
rect 314 -200 372 -188
rect 412 188 470 200
rect 412 -188 424 188
rect 458 -188 470 188
rect 412 -200 470 -188
rect 510 188 568 200
rect 510 -188 522 188
rect 556 -188 568 188
rect 510 -200 568 -188
rect 608 188 666 200
rect 608 -188 620 188
rect 654 -188 666 188
rect 608 -200 666 -188
rect 706 188 764 200
rect 706 -188 718 188
rect 752 -188 764 188
rect 706 -200 764 -188
<< ndiffc >>
rect -752 -188 -718 188
rect -654 -188 -620 188
rect -556 -188 -522 188
rect -458 -188 -424 188
rect -360 -188 -326 188
rect -262 -188 -228 188
rect -164 -188 -130 188
rect -66 -188 -32 188
rect 32 -188 66 188
rect 130 -188 164 188
rect 228 -188 262 188
rect 326 -188 360 188
rect 424 -188 458 188
rect 522 -188 556 188
rect 620 -188 654 188
rect 718 -188 752 188
<< psubdiff >>
rect -866 340 -770 374
rect 770 340 866 374
rect -866 278 -832 340
rect 832 278 866 340
rect -866 -340 -832 -278
rect 832 -340 866 -278
rect -866 -374 -770 -340
rect 770 -374 866 -340
<< psubdiffcont >>
rect -770 340 770 374
rect -866 -278 -832 278
rect 832 -278 866 278
rect -770 -374 770 -340
<< poly >>
rect -621 272 -555 288
rect -621 238 -605 272
rect -571 238 -555 272
rect -706 200 -666 226
rect -621 222 -555 238
rect -425 272 -359 288
rect -425 238 -409 272
rect -375 238 -359 272
rect -608 200 -568 222
rect -510 200 -470 226
rect -425 222 -359 238
rect -229 272 -163 288
rect -229 238 -213 272
rect -179 238 -163 272
rect -412 200 -372 222
rect -314 200 -274 226
rect -229 222 -163 238
rect -33 272 33 288
rect -33 238 -17 272
rect 17 238 33 272
rect -216 200 -176 222
rect -118 200 -78 226
rect -33 222 33 238
rect 163 272 229 288
rect 163 238 179 272
rect 213 238 229 272
rect -20 200 20 222
rect 78 200 118 226
rect 163 222 229 238
rect 359 272 425 288
rect 359 238 375 272
rect 409 238 425 272
rect 176 200 216 222
rect 274 200 314 226
rect 359 222 425 238
rect 555 272 621 288
rect 555 238 571 272
rect 605 238 621 272
rect 372 200 412 222
rect 470 200 510 226
rect 555 222 621 238
rect 568 200 608 222
rect 666 200 706 226
rect -706 -222 -666 -200
rect -719 -238 -653 -222
rect -608 -226 -568 -200
rect -510 -222 -470 -200
rect -719 -272 -703 -238
rect -669 -272 -653 -238
rect -719 -288 -653 -272
rect -523 -238 -457 -222
rect -412 -226 -372 -200
rect -314 -222 -274 -200
rect -523 -272 -507 -238
rect -473 -272 -457 -238
rect -523 -288 -457 -272
rect -327 -238 -261 -222
rect -216 -226 -176 -200
rect -118 -222 -78 -200
rect -327 -272 -311 -238
rect -277 -272 -261 -238
rect -327 -288 -261 -272
rect -131 -238 -65 -222
rect -20 -226 20 -200
rect 78 -222 118 -200
rect -131 -272 -115 -238
rect -81 -272 -65 -238
rect -131 -288 -65 -272
rect 65 -238 131 -222
rect 176 -226 216 -200
rect 274 -222 314 -200
rect 65 -272 81 -238
rect 115 -272 131 -238
rect 65 -288 131 -272
rect 261 -238 327 -222
rect 372 -226 412 -200
rect 470 -222 510 -200
rect 261 -272 277 -238
rect 311 -272 327 -238
rect 261 -288 327 -272
rect 457 -238 523 -222
rect 568 -226 608 -200
rect 666 -222 706 -200
rect 457 -272 473 -238
rect 507 -272 523 -238
rect 457 -288 523 -272
rect 653 -238 719 -222
rect 653 -272 669 -238
rect 703 -272 719 -238
rect 653 -288 719 -272
<< polycont >>
rect -605 238 -571 272
rect -409 238 -375 272
rect -213 238 -179 272
rect -17 238 17 272
rect 179 238 213 272
rect 375 238 409 272
rect 571 238 605 272
rect -703 -272 -669 -238
rect -507 -272 -473 -238
rect -311 -272 -277 -238
rect -115 -272 -81 -238
rect 81 -272 115 -238
rect 277 -272 311 -238
rect 473 -272 507 -238
rect 669 -272 703 -238
<< locali >>
rect -866 340 -770 374
rect 770 340 866 374
rect -866 278 -832 340
rect 832 278 866 340
rect -621 238 -605 272
rect -571 238 -555 272
rect -425 238 -409 272
rect -375 238 -359 272
rect -229 238 -213 272
rect -179 238 -163 272
rect -33 238 -17 272
rect 17 238 33 272
rect 163 238 179 272
rect 213 238 229 272
rect 359 238 375 272
rect 409 238 425 272
rect 555 238 571 272
rect 605 238 621 272
rect -752 188 -718 204
rect -752 -204 -718 -188
rect -654 188 -620 204
rect -654 -204 -620 -188
rect -556 188 -522 204
rect -556 -204 -522 -188
rect -458 188 -424 204
rect -458 -204 -424 -188
rect -360 188 -326 204
rect -360 -204 -326 -188
rect -262 188 -228 204
rect -262 -204 -228 -188
rect -164 188 -130 204
rect -164 -204 -130 -188
rect -66 188 -32 204
rect -66 -204 -32 -188
rect 32 188 66 204
rect 32 -204 66 -188
rect 130 188 164 204
rect 130 -204 164 -188
rect 228 188 262 204
rect 228 -204 262 -188
rect 326 188 360 204
rect 326 -204 360 -188
rect 424 188 458 204
rect 424 -204 458 -188
rect 522 188 556 204
rect 522 -204 556 -188
rect 620 188 654 204
rect 620 -204 654 -188
rect 718 188 752 204
rect 718 -204 752 -188
rect -719 -272 -703 -238
rect -669 -272 -653 -238
rect -523 -272 -507 -238
rect -473 -272 -457 -238
rect -327 -272 -311 -238
rect -277 -272 -261 -238
rect -131 -272 -115 -238
rect -81 -272 -65 -238
rect 65 -272 81 -238
rect 115 -272 131 -238
rect 261 -272 277 -238
rect 311 -272 327 -238
rect 457 -272 473 -238
rect 507 -272 523 -238
rect 653 -272 669 -238
rect 703 -272 719 -238
rect -866 -340 -832 -278
rect 832 -340 866 -278
rect -866 -374 -770 -340
rect 770 -374 866 -340
<< viali >>
rect -605 238 -571 272
rect -409 238 -375 272
rect -213 238 -179 272
rect -17 238 17 272
rect 179 238 213 272
rect 375 238 409 272
rect 571 238 605 272
rect -752 -188 -718 188
rect -654 -188 -620 188
rect -556 -188 -522 188
rect -458 -188 -424 188
rect -360 -188 -326 188
rect -262 -188 -228 188
rect -164 -188 -130 188
rect -66 -188 -32 188
rect 32 -188 66 188
rect 130 -188 164 188
rect 228 -188 262 188
rect 326 -188 360 188
rect 424 -188 458 188
rect 522 -188 556 188
rect 620 -188 654 188
rect 718 -188 752 188
rect -703 -272 -669 -238
rect -507 -272 -473 -238
rect -311 -272 -277 -238
rect -115 -272 -81 -238
rect 81 -272 115 -238
rect 277 -272 311 -238
rect 473 -272 507 -238
rect 669 -272 703 -238
<< metal1 >>
rect -617 272 -559 278
rect -617 238 -605 272
rect -571 238 -559 272
rect -617 232 -559 238
rect -421 272 -363 278
rect -421 238 -409 272
rect -375 238 -363 272
rect -421 232 -363 238
rect -225 272 -167 278
rect -225 238 -213 272
rect -179 238 -167 272
rect -225 232 -167 238
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect 167 272 225 278
rect 167 238 179 272
rect 213 238 225 272
rect 167 232 225 238
rect 363 272 421 278
rect 363 238 375 272
rect 409 238 421 272
rect 363 232 421 238
rect 559 272 617 278
rect 559 238 571 272
rect 605 238 617 272
rect 559 232 617 238
rect -758 188 -712 200
rect -758 -188 -752 188
rect -718 -188 -712 188
rect -758 -200 -712 -188
rect -660 188 -614 200
rect -660 -188 -654 188
rect -620 -188 -614 188
rect -660 -200 -614 -188
rect -562 188 -516 200
rect -562 -188 -556 188
rect -522 -188 -516 188
rect -562 -200 -516 -188
rect -464 188 -418 200
rect -464 -188 -458 188
rect -424 -188 -418 188
rect -464 -200 -418 -188
rect -366 188 -320 200
rect -366 -188 -360 188
rect -326 -188 -320 188
rect -366 -200 -320 -188
rect -268 188 -222 200
rect -268 -188 -262 188
rect -228 -188 -222 188
rect -268 -200 -222 -188
rect -170 188 -124 200
rect -170 -188 -164 188
rect -130 -188 -124 188
rect -170 -200 -124 -188
rect -72 188 -26 200
rect -72 -188 -66 188
rect -32 -188 -26 188
rect -72 -200 -26 -188
rect 26 188 72 200
rect 26 -188 32 188
rect 66 -188 72 188
rect 26 -200 72 -188
rect 124 188 170 200
rect 124 -188 130 188
rect 164 -188 170 188
rect 124 -200 170 -188
rect 222 188 268 200
rect 222 -188 228 188
rect 262 -188 268 188
rect 222 -200 268 -188
rect 320 188 366 200
rect 320 -188 326 188
rect 360 -188 366 188
rect 320 -200 366 -188
rect 418 188 464 200
rect 418 -188 424 188
rect 458 -188 464 188
rect 418 -200 464 -188
rect 516 188 562 200
rect 516 -188 522 188
rect 556 -188 562 188
rect 516 -200 562 -188
rect 614 188 660 200
rect 614 -188 620 188
rect 654 -188 660 188
rect 614 -200 660 -188
rect 712 188 758 200
rect 712 -188 718 188
rect 752 -188 758 188
rect 712 -200 758 -188
rect -715 -238 -657 -232
rect -715 -272 -703 -238
rect -669 -272 -657 -238
rect -715 -278 -657 -272
rect -519 -238 -461 -232
rect -519 -272 -507 -238
rect -473 -272 -461 -238
rect -519 -278 -461 -272
rect -323 -238 -265 -232
rect -323 -272 -311 -238
rect -277 -272 -265 -238
rect -323 -278 -265 -272
rect -127 -238 -69 -232
rect -127 -272 -115 -238
rect -81 -272 -69 -238
rect -127 -278 -69 -272
rect 69 -238 127 -232
rect 69 -272 81 -238
rect 115 -272 127 -238
rect 69 -278 127 -272
rect 265 -238 323 -232
rect 265 -272 277 -238
rect 311 -272 323 -238
rect 265 -278 323 -272
rect 461 -238 519 -232
rect 461 -272 473 -238
rect 507 -272 519 -238
rect 461 -278 519 -272
rect 657 -238 715 -232
rect 657 -272 669 -238
rect 703 -272 715 -238
rect 657 -278 715 -272
<< properties >>
string FIXED_BBOX -849 -357 849 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.2 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
