magic
tech sky130A
magscale 1 2
timestamp 1647868710
<< metal3 >>
rect -1650 1272 1649 1300
rect -1650 -1272 1565 1272
rect 1629 -1272 1649 1272
rect -1650 -1300 1649 -1272
<< via3 >>
rect 1565 -1272 1629 1272
<< mimcap >>
rect -1550 1160 1450 1200
rect -1550 -1160 -1510 1160
rect 1410 -1160 1450 1160
rect -1550 -1200 1450 -1160
<< mimcapcontact >>
rect -1510 -1160 1410 1160
<< metal4 >>
rect 1549 1272 1645 1288
rect -1511 1160 1411 1161
rect -1511 -1160 -1510 1160
rect 1410 -1160 1411 1160
rect -1511 -1161 1411 -1160
rect 1549 -1272 1565 1272
rect 1629 -1272 1645 1272
rect 1549 -1288 1645 -1272
<< properties >>
string FIXED_BBOX -1650 -1300 1550 1300
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15 l 12 val 370.26 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
