magic
tech sky130A
timestamp 1645462850
<< pwell >>
rect -398 -305 398 305
<< nmos >>
rect -300 -200 300 200
<< ndiff >>
rect -329 194 -300 200
rect -329 -194 -323 194
rect -306 -194 -300 194
rect -329 -200 -300 -194
rect 300 194 329 200
rect 300 -194 306 194
rect 323 -194 329 194
rect 300 -200 329 -194
<< ndiffc >>
rect -323 -194 -306 194
rect 306 -194 323 194
<< psubdiff >>
rect -380 270 -332 287
rect 332 270 380 287
rect -380 239 -363 270
rect 363 239 380 270
rect -380 -270 -363 -239
rect 363 -270 380 -239
rect -380 -287 -332 -270
rect 332 -287 380 -270
<< psubdiffcont >>
rect -332 270 332 287
rect -380 -239 -363 239
rect 363 -239 380 239
rect -332 -287 332 -270
<< poly >>
rect -300 236 300 244
rect -300 219 -292 236
rect 292 219 300 236
rect -300 200 300 219
rect -300 -219 300 -200
rect -300 -236 -292 -219
rect 292 -236 300 -219
rect -300 -244 300 -236
<< polycont >>
rect -292 219 292 236
rect -292 -236 292 -219
<< locali >>
rect -380 270 -332 287
rect 332 270 380 287
rect -380 239 -363 270
rect 363 239 380 270
rect -300 219 -292 236
rect 292 219 300 236
rect -323 194 -306 202
rect -323 -202 -306 -194
rect 306 194 323 202
rect 306 -202 323 -194
rect -300 -236 -292 -219
rect 292 -236 300 -219
rect -380 -270 -363 -239
rect 363 -270 380 -239
rect -380 -287 -332 -270
rect 332 -287 380 -270
<< viali >>
rect -292 219 292 236
rect -323 -194 -306 194
rect 306 -194 323 194
rect -292 -236 292 -219
<< metal1 >>
rect -298 236 298 239
rect -298 219 -292 236
rect 292 219 298 236
rect -298 216 298 219
rect -326 194 -303 200
rect -326 -194 -323 194
rect -306 -194 -303 194
rect -326 -200 -303 -194
rect 303 194 326 200
rect 303 -194 306 194
rect 323 -194 326 194
rect 303 -200 326 -194
rect -298 -219 298 -216
rect -298 -236 -292 -219
rect 292 -236 298 -219
rect -298 -239 298 -236
<< properties >>
string FIXED_BBOX -371 -278 371 278
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
