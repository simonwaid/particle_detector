magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< pwell >>
rect 32 2696 1154 2762
rect 32 2186 1154 2252
rect 32 2078 1154 2144
rect 86 1906 1100 2066
rect 32 1568 1154 1634
rect 32 1460 1154 1526
rect 32 950 1154 1016
rect 32 842 1154 908
rect 32 332 1154 398
rect 42 42 1410 88
rect 42 -468 1408 -422
<< poly >>
rect 32 2746 1154 2762
rect 32 2712 144 2746
rect 178 2712 336 2746
rect 370 2712 528 2746
rect 562 2712 720 2746
rect 754 2712 912 2746
rect 946 2712 1104 2746
rect 1138 2712 1154 2746
rect 32 2696 1154 2712
rect 32 2236 1154 2252
rect 32 2202 48 2236
rect 82 2202 240 2236
rect 274 2202 432 2236
rect 466 2202 624 2236
rect 658 2202 816 2236
rect 850 2202 1008 2236
rect 1042 2202 1154 2236
rect 32 2186 1154 2202
rect 32 2128 1154 2144
rect 32 2094 48 2128
rect 82 2094 240 2128
rect 274 2094 432 2128
rect 466 2094 624 2128
rect 658 2094 816 2128
rect 850 2094 1008 2128
rect 1042 2094 1154 2128
rect 32 2078 1154 2094
rect 32 1618 1154 1634
rect 32 1584 144 1618
rect 178 1584 336 1618
rect 370 1584 528 1618
rect 562 1584 720 1618
rect 754 1584 912 1618
rect 946 1584 1104 1618
rect 1138 1584 1154 1618
rect 32 1568 1154 1584
rect 32 1510 1154 1526
rect 32 1476 144 1510
rect 178 1476 336 1510
rect 370 1476 528 1510
rect 562 1476 720 1510
rect 754 1476 912 1510
rect 946 1476 1104 1510
rect 1138 1476 1154 1510
rect 32 1460 1154 1476
rect 32 1000 1154 1016
rect 32 966 48 1000
rect 82 966 240 1000
rect 274 966 432 1000
rect 466 966 624 1000
rect 658 966 816 1000
rect 850 966 1008 1000
rect 1042 966 1154 1000
rect 32 950 1154 966
rect 32 892 1154 908
rect 32 858 48 892
rect 82 858 240 892
rect 274 858 432 892
rect 466 858 624 892
rect 658 858 816 892
rect 850 858 1008 892
rect 1042 858 1154 892
rect 32 842 1154 858
rect 32 382 1154 398
rect 32 348 144 382
rect 178 348 336 382
rect 370 348 528 382
rect 562 348 720 382
rect 754 348 912 382
rect 946 348 1104 382
rect 1138 348 1154 382
rect 32 332 1154 348
rect 42 42 1410 88
rect 42 -468 1408 -422
<< polycont >>
rect 144 2712 178 2746
rect 336 2712 370 2746
rect 528 2712 562 2746
rect 720 2712 754 2746
rect 912 2712 946 2746
rect 1104 2712 1138 2746
rect 48 2202 82 2236
rect 240 2202 274 2236
rect 432 2202 466 2236
rect 624 2202 658 2236
rect 816 2202 850 2236
rect 1008 2202 1042 2236
rect 48 2094 82 2128
rect 240 2094 274 2128
rect 432 2094 466 2128
rect 624 2094 658 2128
rect 816 2094 850 2128
rect 1008 2094 1042 2128
rect 144 1584 178 1618
rect 336 1584 370 1618
rect 528 1584 562 1618
rect 720 1584 754 1618
rect 912 1584 946 1618
rect 1104 1584 1138 1618
rect 144 1476 178 1510
rect 336 1476 370 1510
rect 528 1476 562 1510
rect 720 1476 754 1510
rect 912 1476 946 1510
rect 1104 1476 1138 1510
rect 48 966 82 1000
rect 240 966 274 1000
rect 432 966 466 1000
rect 624 966 658 1000
rect 816 966 850 1000
rect 1008 966 1042 1000
rect 48 858 82 892
rect 240 858 274 892
rect 432 858 466 892
rect 624 858 658 892
rect 816 858 850 892
rect 1008 858 1042 892
rect 144 348 178 382
rect 336 348 370 382
rect 528 348 562 382
rect 720 348 754 382
rect 912 348 946 382
rect 1104 348 1138 382
<< locali >>
rect 32 2712 144 2746
rect 178 2712 336 2746
rect 370 2712 528 2746
rect 562 2712 720 2746
rect 754 2712 912 2746
rect 946 2712 1104 2746
rect 1138 2712 1154 2746
rect 32 2202 48 2236
rect 82 2202 240 2236
rect 274 2202 432 2236
rect 466 2202 624 2236
rect 658 2202 816 2236
rect 850 2202 1008 2236
rect 1042 2202 1154 2236
rect 32 2094 48 2128
rect 82 2094 240 2128
rect 274 2094 432 2128
rect 466 2094 624 2128
rect 658 2094 816 2128
rect 850 2094 1008 2128
rect 1042 2094 1154 2128
rect 32 1584 144 1618
rect 178 1584 336 1618
rect 370 1584 528 1618
rect 562 1584 720 1618
rect 754 1584 912 1618
rect 946 1584 1104 1618
rect 1138 1584 1154 1618
rect 32 1476 144 1510
rect 178 1476 336 1510
rect 370 1476 528 1510
rect 562 1476 720 1510
rect 754 1476 912 1510
rect 946 1476 1104 1510
rect 1138 1476 1154 1510
rect 32 966 48 1000
rect 82 966 240 1000
rect 274 966 432 1000
rect 466 966 624 1000
rect 658 966 816 1000
rect 850 966 1008 1000
rect 1042 966 1154 1000
rect 32 858 48 892
rect 82 858 240 892
rect 274 858 432 892
rect 466 858 624 892
rect 658 858 816 892
rect 850 858 1008 892
rect 1042 858 1154 892
rect 32 348 144 382
rect 178 348 336 382
rect 370 348 528 382
rect 562 348 720 382
rect 754 348 912 382
rect 946 348 1104 382
rect 1138 348 1154 382
rect 1290 260 1520 2840
rect -110 170 1520 260
rect -100 10 -60 170
rect 1290 160 1520 170
rect 42 48 1408 82
rect 1500 10 1550 160
rect -100 -390 10 10
rect 1450 -390 1550 10
rect 42 -462 1408 -428
<< viali >>
rect 144 2712 178 2746
rect 336 2712 370 2746
rect 528 2712 562 2746
rect 720 2712 754 2746
rect 912 2712 946 2746
rect 1104 2712 1138 2746
rect 48 2202 82 2236
rect 240 2202 274 2236
rect 432 2202 466 2236
rect 624 2202 658 2236
rect 816 2202 850 2236
rect 1008 2202 1042 2236
rect 48 2094 82 2128
rect 240 2094 274 2128
rect 432 2094 466 2128
rect 624 2094 658 2128
rect 816 2094 850 2128
rect 1008 2094 1042 2128
rect 144 1584 178 1618
rect 336 1584 370 1618
rect 528 1584 562 1618
rect 720 1584 754 1618
rect 912 1584 946 1618
rect 1104 1584 1138 1618
rect 144 1476 178 1510
rect 336 1476 370 1510
rect 528 1476 562 1510
rect 720 1476 754 1510
rect 912 1476 946 1510
rect 1104 1476 1138 1510
rect 48 966 82 1000
rect 240 966 274 1000
rect 432 966 466 1000
rect 624 966 658 1000
rect 816 966 850 1000
rect 1008 966 1042 1000
rect 48 858 82 892
rect 240 858 274 892
rect 432 858 466 892
rect 624 858 658 892
rect 816 858 850 892
rect 1008 858 1042 892
rect 144 348 178 382
rect 336 348 370 382
rect 528 348 562 382
rect 720 348 754 382
rect 912 348 946 382
rect 1104 348 1138 382
rect -10 -580 160 -510
rect 1280 -580 1450 -510
<< metal1 >>
rect -120 2746 1310 2760
rect -120 2712 144 2746
rect 178 2712 336 2746
rect 370 2712 528 2746
rect 562 2712 720 2746
rect 754 2712 912 2746
rect 946 2712 1104 2746
rect 1138 2712 1310 2746
rect -120 2710 1310 2712
rect -120 2240 -50 2710
rect 32 2706 1154 2710
rect 76 2498 86 2674
rect 140 2498 150 2674
rect 268 2498 278 2674
rect 332 2498 342 2674
rect 460 2498 470 2674
rect 524 2498 534 2674
rect 652 2498 662 2674
rect 716 2498 726 2674
rect 844 2498 854 2674
rect 908 2498 918 2674
rect 1036 2498 1046 2674
rect 1100 2498 1110 2674
rect -20 2274 -10 2450
rect 44 2274 54 2450
rect 172 2274 182 2450
rect 236 2274 246 2450
rect 364 2274 374 2450
rect 428 2274 438 2450
rect 556 2274 566 2450
rect 620 2274 630 2450
rect 748 2274 758 2450
rect 812 2274 822 2450
rect 940 2274 950 2450
rect 1004 2274 1014 2450
rect 1132 2274 1142 2450
rect 1196 2274 1206 2450
rect 32 2240 1154 2242
rect 1240 2240 1310 2710
rect -120 2236 1310 2240
rect -120 2202 48 2236
rect 82 2202 240 2236
rect 274 2202 432 2236
rect 466 2202 624 2236
rect 658 2202 816 2236
rect 850 2202 1008 2236
rect 1042 2202 1310 2236
rect -120 2190 1310 2202
rect -120 2140 -50 2190
rect 1240 2140 1310 2190
rect -120 2128 1310 2140
rect -120 2094 48 2128
rect 82 2094 240 2128
rect 274 2094 432 2128
rect 466 2094 624 2128
rect 658 2094 816 2128
rect 850 2094 1008 2128
rect 1042 2094 1310 2128
rect -120 2090 1310 2094
rect -120 1620 -50 2090
rect 32 2088 1154 2090
rect 76 1880 86 2056
rect 140 1880 150 2056
rect 268 1880 278 2056
rect 332 1880 342 2056
rect 460 1880 470 2056
rect 524 1880 534 2056
rect 652 1880 662 2056
rect 716 1880 726 2056
rect 844 1880 854 2056
rect 908 1880 918 2056
rect 1036 1880 1046 2056
rect 1100 1880 1110 2056
rect -20 1656 -10 1832
rect 44 1656 54 1832
rect 172 1656 182 1832
rect 236 1656 246 1832
rect 364 1656 374 1832
rect 428 1656 438 1832
rect 556 1656 566 1832
rect 620 1656 630 1832
rect 748 1656 758 1832
rect 812 1656 822 1832
rect 940 1656 950 1832
rect 1004 1656 1014 1832
rect 1132 1656 1142 1832
rect 1196 1656 1206 1832
rect 32 1620 1154 1624
rect 1240 1620 1310 2090
rect -120 1618 1310 1620
rect -120 1584 144 1618
rect 178 1584 336 1618
rect 370 1584 528 1618
rect 562 1584 720 1618
rect 754 1584 912 1618
rect 946 1584 1104 1618
rect 1138 1584 1310 1618
rect -120 1570 1310 1584
rect -120 1520 -50 1570
rect 1240 1520 1310 1570
rect -120 1510 1310 1520
rect -120 1476 144 1510
rect 178 1476 336 1510
rect 370 1476 528 1510
rect 562 1476 720 1510
rect 754 1476 912 1510
rect 946 1476 1104 1510
rect 1138 1476 1310 1510
rect -120 1470 1310 1476
rect -120 1010 -50 1470
rect 76 1262 86 1438
rect 140 1262 150 1438
rect 268 1262 278 1438
rect 332 1262 342 1438
rect 460 1262 470 1438
rect 524 1262 534 1438
rect 652 1262 662 1438
rect 716 1262 726 1438
rect 844 1262 854 1438
rect 908 1262 918 1438
rect 1036 1262 1046 1438
rect 1100 1262 1110 1438
rect -20 1038 -10 1214
rect 44 1038 54 1214
rect 172 1038 182 1214
rect 236 1038 246 1214
rect 364 1038 374 1214
rect 428 1038 438 1214
rect 556 1038 566 1214
rect 620 1038 630 1214
rect 748 1038 758 1214
rect 812 1038 822 1214
rect 940 1038 950 1214
rect 1004 1038 1014 1214
rect 1132 1038 1142 1214
rect 1196 1038 1206 1214
rect 1240 1010 1310 1470
rect -120 1000 1310 1010
rect -120 966 48 1000
rect 82 966 240 1000
rect 274 966 432 1000
rect 466 966 624 1000
rect 658 966 816 1000
rect 850 966 1008 1000
rect 1042 966 1310 1000
rect -120 960 1310 966
rect -120 900 -50 960
rect 1240 900 1310 960
rect -120 892 1310 900
rect -120 858 48 892
rect 82 858 240 892
rect 274 858 432 892
rect 466 858 624 892
rect 658 858 816 892
rect 850 858 1008 892
rect 1042 858 1310 892
rect -120 850 1310 858
rect -120 390 -50 850
rect 76 644 86 820
rect 140 644 150 820
rect 268 644 278 820
rect 332 644 342 820
rect 460 644 470 820
rect 524 644 534 820
rect 652 644 662 820
rect 716 644 726 820
rect 844 644 854 820
rect 908 644 918 820
rect 1036 644 1046 820
rect 1100 644 1110 820
rect -20 420 -10 596
rect 44 420 54 596
rect 172 420 182 596
rect 236 420 246 596
rect 364 420 374 596
rect 428 420 438 596
rect 556 420 566 596
rect 620 420 630 596
rect 748 420 758 596
rect 812 420 822 596
rect 940 420 950 596
rect 1004 420 1014 596
rect 1132 420 1142 596
rect 1196 420 1206 596
rect 1240 390 1310 850
rect -120 382 1310 390
rect -120 348 144 382
rect 178 348 336 382
rect 370 348 528 382
rect 562 348 720 382
rect 754 348 912 382
rect 946 348 1104 382
rect 1138 348 1310 382
rect -120 340 1310 348
rect -120 90 -50 340
rect 1240 90 1310 340
rect -120 40 1570 90
rect -120 -420 -50 40
rect 98 -166 108 10
rect 162 -166 172 10
rect 334 -166 344 10
rect 398 -166 408 10
rect 570 -166 580 10
rect 634 -166 644 10
rect 806 -166 816 10
rect 870 -166 880 10
rect 1042 -166 1052 10
rect 1106 -166 1116 10
rect 1278 -166 1288 10
rect 1342 -166 1352 10
rect -20 -390 -10 -214
rect 44 -390 54 -214
rect 216 -390 226 -214
rect 280 -390 290 -214
rect 452 -390 462 -214
rect 516 -390 526 -214
rect 688 -390 698 -214
rect 752 -390 762 -214
rect 924 -390 934 -214
rect 988 -390 998 -214
rect 1160 -390 1170 -214
rect 1224 -390 1234 -214
rect 1396 -390 1406 -214
rect 1460 -390 1470 -214
rect 1500 -420 1570 40
rect -120 -470 1570 -420
rect -22 -510 172 -504
rect -22 -580 -10 -510
rect 160 -580 172 -510
rect -22 -586 172 -580
rect 1268 -510 1462 -504
rect 1268 -580 1280 -510
rect 1450 -580 1462 -510
rect 1268 -586 1462 -580
<< via1 >>
rect 86 2498 140 2674
rect 278 2498 332 2674
rect 470 2498 524 2674
rect 662 2498 716 2674
rect 854 2498 908 2674
rect 1046 2498 1100 2674
rect -10 2274 44 2450
rect 182 2274 236 2450
rect 374 2274 428 2450
rect 566 2274 620 2450
rect 758 2274 812 2450
rect 950 2274 1004 2450
rect 1142 2274 1196 2450
rect 86 1880 140 2056
rect 278 1880 332 2056
rect 470 1880 524 2056
rect 662 1880 716 2056
rect 854 1880 908 2056
rect 1046 1880 1100 2056
rect -10 1656 44 1832
rect 182 1656 236 1832
rect 374 1656 428 1832
rect 566 1656 620 1832
rect 758 1656 812 1832
rect 950 1656 1004 1832
rect 1142 1656 1196 1832
rect 86 1262 140 1438
rect 278 1262 332 1438
rect 470 1262 524 1438
rect 662 1262 716 1438
rect 854 1262 908 1438
rect 1046 1262 1100 1438
rect -10 1038 44 1214
rect 182 1038 236 1214
rect 374 1038 428 1214
rect 566 1038 620 1214
rect 758 1038 812 1214
rect 950 1038 1004 1214
rect 1142 1038 1196 1214
rect 86 644 140 820
rect 278 644 332 820
rect 470 644 524 820
rect 662 644 716 820
rect 854 644 908 820
rect 1046 644 1100 820
rect -10 420 44 596
rect 182 420 236 596
rect 374 420 428 596
rect 566 420 620 596
rect 758 420 812 596
rect 950 420 1004 596
rect 1142 420 1196 596
rect 108 -166 162 10
rect 344 -166 398 10
rect 580 -166 634 10
rect 816 -166 870 10
rect 1052 -166 1106 10
rect 1288 -166 1342 10
rect -10 -390 44 -214
rect 226 -390 280 -214
rect 462 -390 516 -214
rect 698 -390 752 -214
rect 934 -390 988 -214
rect 1170 -390 1224 -214
rect 1406 -390 1460 -214
rect -10 -580 160 -510
rect 1280 -580 1450 -510
<< metal2 >>
rect -70 2700 1100 2740
rect 620 2674 1100 2700
rect 620 2540 662 2674
rect -70 2520 86 2540
rect 140 2520 278 2540
rect 86 2488 140 2498
rect 332 2520 470 2540
rect 278 2488 332 2498
rect 524 2520 662 2540
rect 470 2488 524 2498
rect 716 2520 854 2674
rect 662 2488 716 2498
rect 908 2520 1046 2674
rect 854 2488 908 2498
rect 1046 2488 1100 2498
rect -10 2450 44 2460
rect 182 2450 236 2460
rect 44 2274 182 2424
rect 374 2450 428 2460
rect 236 2274 374 2424
rect 566 2450 620 2460
rect 428 2274 566 2424
rect 758 2450 812 2460
rect 730 2424 758 2430
rect 620 2420 758 2424
rect 950 2450 1004 2460
rect 812 2420 950 2430
rect 1142 2450 1196 2460
rect 1004 2420 1142 2430
rect 1196 2420 1460 2430
rect 620 2274 730 2420
rect -10 2260 730 2274
rect -10 2170 1460 2260
rect -70 2080 1100 2130
rect 620 2056 1100 2080
rect 620 1920 662 2056
rect -70 1910 86 1920
rect 140 1906 278 1920
rect 86 1870 140 1880
rect 332 1906 470 1920
rect 278 1870 332 1880
rect 524 1906 662 1920
rect 470 1870 524 1880
rect 716 1906 854 2056
rect 662 1870 716 1880
rect 908 1906 1046 2056
rect 854 1870 908 1880
rect 1046 1870 1100 1880
rect -10 1832 44 1842
rect 182 1832 236 1842
rect 44 1656 182 1810
rect 374 1832 428 1842
rect 236 1656 374 1810
rect 566 1832 620 1842
rect 428 1656 566 1810
rect 758 1832 812 1842
rect 620 1800 758 1810
rect 950 1832 1004 1842
rect 812 1800 950 1810
rect 1142 1832 1196 1842
rect 1004 1800 1142 1810
rect 1196 1800 1460 1810
rect 620 1656 730 1800
rect -10 1640 730 1656
rect -10 1560 1460 1640
rect -70 1460 1100 1510
rect 620 1438 1100 1460
rect 620 1300 662 1438
rect -70 1290 86 1300
rect 140 1288 278 1300
rect 86 1252 140 1262
rect 332 1288 470 1300
rect 278 1252 332 1262
rect 524 1288 662 1300
rect 470 1252 524 1262
rect 716 1288 854 1438
rect 662 1252 716 1262
rect 908 1288 1046 1438
rect 854 1252 908 1262
rect 1046 1252 1100 1262
rect -10 1214 44 1224
rect 182 1214 236 1224
rect 44 1038 182 1190
rect 374 1214 428 1224
rect 236 1038 374 1190
rect 566 1214 620 1224
rect 428 1038 566 1190
rect 758 1214 812 1224
rect 620 1180 758 1190
rect 950 1214 1004 1224
rect 812 1180 950 1190
rect 1142 1214 1196 1224
rect 1004 1180 1142 1190
rect 1196 1180 1460 1190
rect 620 1038 730 1180
rect -10 1020 730 1038
rect -10 940 1460 1020
rect -70 840 1100 890
rect 620 820 1100 840
rect 620 680 662 820
rect -70 670 86 680
rect 140 670 278 680
rect 86 634 140 644
rect 332 670 470 680
rect 278 634 332 644
rect 524 670 662 680
rect 470 634 524 644
rect 716 670 854 820
rect 662 634 716 644
rect 908 670 1046 820
rect 854 634 908 644
rect 1046 634 1100 644
rect -10 596 44 606
rect 182 596 236 606
rect 44 420 182 570
rect 374 596 428 606
rect 236 420 374 570
rect 566 596 620 606
rect 428 420 566 570
rect 758 596 812 606
rect 620 560 758 570
rect 950 596 1004 606
rect 812 560 950 570
rect 1142 596 1196 606
rect 1004 560 1142 570
rect 1196 560 1460 570
rect 620 420 730 560
rect -10 130 730 420
rect -10 10 1460 130
rect -10 -140 108 10
rect 162 -140 344 10
rect 108 -176 162 -166
rect 398 -140 580 10
rect 344 -176 398 -166
rect 634 -140 816 10
rect 810 -150 816 -140
rect 580 -176 634 -166
rect 870 -140 1052 10
rect 870 -150 880 -140
rect 1040 -150 1052 -140
rect 816 -176 870 -166
rect 1106 -140 1288 10
rect 1106 -150 1120 -140
rect 1280 -150 1288 -140
rect 1052 -176 1106 -166
rect 1342 -140 1460 10
rect 1342 -150 1360 -140
rect 1288 -176 1342 -166
rect -10 -214 44 -204
rect 226 -214 280 -204
rect 44 -390 226 -240
rect 462 -214 516 -204
rect 280 -390 462 -240
rect 698 -214 752 -204
rect 516 -390 698 -240
rect 934 -214 988 -204
rect 752 -390 934 -240
rect 1170 -214 1224 -204
rect 988 -390 1170 -240
rect 1406 -214 1460 -204
rect 1224 -390 1406 -240
rect -10 -400 1460 -390
rect -10 -510 160 -400
rect -10 -590 160 -580
rect 1280 -510 1450 -400
rect 1280 -590 1450 -580
<< via2 >>
rect -70 2674 620 2700
rect -70 2540 86 2674
rect 86 2540 140 2674
rect 140 2540 278 2674
rect 278 2540 332 2674
rect 332 2540 470 2674
rect 470 2540 524 2674
rect 524 2540 620 2674
rect 730 2274 758 2420
rect 758 2274 812 2420
rect 812 2274 950 2420
rect 950 2274 1004 2420
rect 1004 2274 1142 2420
rect 1142 2274 1196 2420
rect 1196 2274 1460 2420
rect 730 2260 1460 2274
rect -70 2056 620 2080
rect -70 1920 86 2056
rect 86 1920 140 2056
rect 140 1920 278 2056
rect 278 1920 332 2056
rect 332 1920 470 2056
rect 470 1920 524 2056
rect 524 1920 620 2056
rect 730 1656 758 1800
rect 758 1656 812 1800
rect 812 1656 950 1800
rect 950 1656 1004 1800
rect 1004 1656 1142 1800
rect 1142 1656 1196 1800
rect 1196 1656 1460 1800
rect 730 1640 1460 1656
rect -70 1438 620 1460
rect -70 1300 86 1438
rect 86 1300 140 1438
rect 140 1300 278 1438
rect 278 1300 332 1438
rect 332 1300 470 1438
rect 470 1300 524 1438
rect 524 1300 620 1438
rect 730 1038 758 1180
rect 758 1038 812 1180
rect 812 1038 950 1180
rect 950 1038 1004 1180
rect 1004 1038 1142 1180
rect 1142 1038 1196 1180
rect 1196 1038 1460 1180
rect 730 1020 1460 1038
rect -70 820 620 840
rect -70 680 86 820
rect 86 680 140 820
rect 140 680 278 820
rect 278 680 332 820
rect 332 680 470 820
rect 470 680 524 820
rect 524 680 620 820
rect 730 420 758 560
rect 758 420 812 560
rect 812 420 950 560
rect 950 420 1004 560
rect 1004 420 1142 560
rect 1142 420 1196 560
rect 1196 420 1460 560
rect 730 130 1460 420
<< metal3 >>
rect -70 2705 620 2710
rect -80 2700 630 2705
rect -80 2540 -70 2700
rect 620 2540 630 2700
rect -80 2535 630 2540
rect -70 2085 620 2535
rect 730 2425 1460 2430
rect 720 2420 1470 2425
rect 720 2260 730 2420
rect 1460 2260 1470 2420
rect 720 2255 1470 2260
rect -80 2080 630 2085
rect -80 1920 -70 2080
rect 620 1920 630 2080
rect -80 1915 630 1920
rect -70 1465 620 1915
rect 730 1805 1460 2255
rect 720 1800 1470 1805
rect 720 1640 730 1800
rect 1460 1640 1470 1800
rect 720 1635 1470 1640
rect -80 1460 630 1465
rect -80 1300 -70 1460
rect 620 1300 630 1460
rect -80 1295 630 1300
rect -70 845 620 1295
rect 730 1185 1460 1635
rect 720 1180 1470 1185
rect 720 1020 730 1180
rect 1460 1020 1470 1180
rect 720 1015 1470 1020
rect -80 840 630 845
rect -80 680 -70 840
rect 620 680 630 840
rect -80 675 630 680
rect -70 670 620 675
rect 730 565 1460 1015
rect 720 560 1470 565
rect 720 130 730 560
rect 1460 130 1470 560
rect 720 125 1470 130
use sky130_fd_pr__nfet_01v8_HR8DH9  sky130_fd_pr__nfet_01v8_HR8DH9_0
timestamp 1654760956
transform 1 0 725 0 1 -190
box -875 -410 875 410
use sky130_fd_pr__nfet_01v8_XZXALN  sky130_fd_pr__nfet_01v8_XZXALN_0
timestamp 1654760956
transform 1 0 593 0 1 1547
box -743 -1337 743 1337
<< end >>
