magic
tech sky130B
magscale 1 2
timestamp 1654611687
<< error_p >>
rect -678 265 -620 271
rect -560 265 -502 271
rect -442 265 -384 271
rect -324 265 -266 271
rect -206 265 -148 271
rect -88 265 -30 271
rect 30 265 88 271
rect 148 265 206 271
rect 266 265 324 271
rect 384 265 442 271
rect 502 265 560 271
rect 620 265 678 271
rect -678 231 -666 265
rect -560 231 -548 265
rect -442 231 -430 265
rect -324 231 -312 265
rect -206 231 -194 265
rect -88 231 -76 265
rect 30 231 42 265
rect 148 231 160 265
rect 266 231 278 265
rect 384 231 396 265
rect 502 231 514 265
rect 620 231 632 265
rect -678 225 -620 231
rect -560 225 -502 231
rect -442 225 -384 231
rect -324 225 -266 231
rect -206 225 -148 231
rect -88 225 -30 231
rect 30 225 88 231
rect 148 225 206 231
rect 266 225 324 231
rect 384 225 442 231
rect 502 225 560 231
rect 620 225 678 231
rect -678 71 -620 77
rect -560 71 -502 77
rect -442 71 -384 77
rect -324 71 -266 77
rect -206 71 -148 77
rect -88 71 -30 77
rect 30 71 88 77
rect 148 71 206 77
rect 266 71 324 77
rect 384 71 442 77
rect 502 71 560 77
rect 620 71 678 77
rect -678 37 -666 71
rect -560 37 -548 71
rect -442 37 -430 71
rect -324 37 -312 71
rect -206 37 -194 71
rect -88 37 -76 71
rect 30 37 42 71
rect 148 37 160 71
rect 266 37 278 71
rect 384 37 396 71
rect 502 37 514 71
rect 620 37 632 71
rect -678 31 -620 37
rect -560 31 -502 37
rect -442 31 -384 37
rect -324 31 -266 37
rect -206 31 -148 37
rect -88 31 -30 37
rect 30 31 88 37
rect 148 31 206 37
rect 266 31 324 37
rect 384 31 442 37
rect 502 31 560 37
rect 620 31 678 37
rect -678 -37 -620 -31
rect -560 -37 -502 -31
rect -442 -37 -384 -31
rect -324 -37 -266 -31
rect -206 -37 -148 -31
rect -88 -37 -30 -31
rect 30 -37 88 -31
rect 148 -37 206 -31
rect 266 -37 324 -31
rect 384 -37 442 -31
rect 502 -37 560 -31
rect 620 -37 678 -31
rect -678 -71 -666 -37
rect -560 -71 -548 -37
rect -442 -71 -430 -37
rect -324 -71 -312 -37
rect -206 -71 -194 -37
rect -88 -71 -76 -37
rect 30 -71 42 -37
rect 148 -71 160 -37
rect 266 -71 278 -37
rect 384 -71 396 -37
rect 502 -71 514 -37
rect 620 -71 632 -37
rect -678 -77 -620 -71
rect -560 -77 -502 -71
rect -442 -77 -384 -71
rect -324 -77 -266 -71
rect -206 -77 -148 -71
rect -88 -77 -30 -71
rect 30 -77 88 -71
rect 148 -77 206 -71
rect 266 -77 324 -71
rect 384 -77 442 -71
rect 502 -77 560 -71
rect 620 -77 678 -71
rect -678 -231 -620 -225
rect -560 -231 -502 -225
rect -442 -231 -384 -225
rect -324 -231 -266 -225
rect -206 -231 -148 -225
rect -88 -231 -30 -225
rect 30 -231 88 -225
rect 148 -231 206 -225
rect 266 -231 324 -225
rect 384 -231 442 -225
rect 502 -231 560 -225
rect 620 -231 678 -225
rect -678 -265 -666 -231
rect -560 -265 -548 -231
rect -442 -265 -430 -231
rect -324 -265 -312 -231
rect -206 -265 -194 -231
rect -88 -265 -76 -231
rect 30 -265 42 -231
rect 148 -265 160 -231
rect 266 -265 278 -231
rect 384 -265 396 -231
rect 502 -265 514 -231
rect 620 -265 632 -231
rect -678 -271 -620 -265
rect -560 -271 -502 -265
rect -442 -271 -384 -265
rect -324 -271 -266 -265
rect -206 -271 -148 -265
rect -88 -271 -30 -265
rect 30 -271 88 -265
rect 148 -271 206 -265
rect 266 -271 324 -265
rect 384 -271 442 -265
rect 502 -271 560 -265
rect 620 -271 678 -265
<< pwell >>
rect -875 -403 875 403
<< nmoslvt >>
rect -679 109 -619 193
rect -561 109 -501 193
rect -443 109 -383 193
rect -325 109 -265 193
rect -207 109 -147 193
rect -89 109 -29 193
rect 29 109 89 193
rect 147 109 207 193
rect 265 109 325 193
rect 383 109 443 193
rect 501 109 561 193
rect 619 109 679 193
rect -679 -193 -619 -109
rect -561 -193 -501 -109
rect -443 -193 -383 -109
rect -325 -193 -265 -109
rect -207 -193 -147 -109
rect -89 -193 -29 -109
rect 29 -193 89 -109
rect 147 -193 207 -109
rect 265 -193 325 -109
rect 383 -193 443 -109
rect 501 -193 561 -109
rect 619 -193 679 -109
<< ndiff >>
rect -737 181 -679 193
rect -737 121 -725 181
rect -691 121 -679 181
rect -737 109 -679 121
rect -619 181 -561 193
rect -619 121 -607 181
rect -573 121 -561 181
rect -619 109 -561 121
rect -501 181 -443 193
rect -501 121 -489 181
rect -455 121 -443 181
rect -501 109 -443 121
rect -383 181 -325 193
rect -383 121 -371 181
rect -337 121 -325 181
rect -383 109 -325 121
rect -265 181 -207 193
rect -265 121 -253 181
rect -219 121 -207 181
rect -265 109 -207 121
rect -147 181 -89 193
rect -147 121 -135 181
rect -101 121 -89 181
rect -147 109 -89 121
rect -29 181 29 193
rect -29 121 -17 181
rect 17 121 29 181
rect -29 109 29 121
rect 89 181 147 193
rect 89 121 101 181
rect 135 121 147 181
rect 89 109 147 121
rect 207 181 265 193
rect 207 121 219 181
rect 253 121 265 181
rect 207 109 265 121
rect 325 181 383 193
rect 325 121 337 181
rect 371 121 383 181
rect 325 109 383 121
rect 443 181 501 193
rect 443 121 455 181
rect 489 121 501 181
rect 443 109 501 121
rect 561 181 619 193
rect 561 121 573 181
rect 607 121 619 181
rect 561 109 619 121
rect 679 181 737 193
rect 679 121 691 181
rect 725 121 737 181
rect 679 109 737 121
rect -737 -121 -679 -109
rect -737 -181 -725 -121
rect -691 -181 -679 -121
rect -737 -193 -679 -181
rect -619 -121 -561 -109
rect -619 -181 -607 -121
rect -573 -181 -561 -121
rect -619 -193 -561 -181
rect -501 -121 -443 -109
rect -501 -181 -489 -121
rect -455 -181 -443 -121
rect -501 -193 -443 -181
rect -383 -121 -325 -109
rect -383 -181 -371 -121
rect -337 -181 -325 -121
rect -383 -193 -325 -181
rect -265 -121 -207 -109
rect -265 -181 -253 -121
rect -219 -181 -207 -121
rect -265 -193 -207 -181
rect -147 -121 -89 -109
rect -147 -181 -135 -121
rect -101 -181 -89 -121
rect -147 -193 -89 -181
rect -29 -121 29 -109
rect -29 -181 -17 -121
rect 17 -181 29 -121
rect -29 -193 29 -181
rect 89 -121 147 -109
rect 89 -181 101 -121
rect 135 -181 147 -121
rect 89 -193 147 -181
rect 207 -121 265 -109
rect 207 -181 219 -121
rect 253 -181 265 -121
rect 207 -193 265 -181
rect 325 -121 383 -109
rect 325 -181 337 -121
rect 371 -181 383 -121
rect 325 -193 383 -181
rect 443 -121 501 -109
rect 443 -181 455 -121
rect 489 -181 501 -121
rect 443 -193 501 -181
rect 561 -121 619 -109
rect 561 -181 573 -121
rect 607 -181 619 -121
rect 561 -193 619 -181
rect 679 -121 737 -109
rect 679 -181 691 -121
rect 725 -181 737 -121
rect 679 -193 737 -181
<< ndiffc >>
rect -725 121 -691 181
rect -607 121 -573 181
rect -489 121 -455 181
rect -371 121 -337 181
rect -253 121 -219 181
rect -135 121 -101 181
rect -17 121 17 181
rect 101 121 135 181
rect 219 121 253 181
rect 337 121 371 181
rect 455 121 489 181
rect 573 121 607 181
rect 691 121 725 181
rect -725 -181 -691 -121
rect -607 -181 -573 -121
rect -489 -181 -455 -121
rect -371 -181 -337 -121
rect -253 -181 -219 -121
rect -135 -181 -101 -121
rect -17 -181 17 -121
rect 101 -181 135 -121
rect 219 -181 253 -121
rect 337 -181 371 -121
rect 455 -181 489 -121
rect 573 -181 607 -121
rect 691 -181 725 -121
<< psubdiff >>
rect -839 333 -743 367
rect 743 333 839 367
rect -839 271 -805 333
rect 805 271 839 333
rect -839 -333 -805 -271
rect 805 -333 839 -271
rect -839 -367 -743 -333
rect 743 -367 839 -333
<< psubdiffcont >>
rect -743 333 743 367
rect -839 -271 -805 271
rect 805 -271 839 271
rect -743 -367 743 -333
<< poly >>
rect -682 265 -616 281
rect -682 231 -666 265
rect -632 231 -616 265
rect -682 215 -616 231
rect -564 265 -498 281
rect -564 231 -548 265
rect -514 231 -498 265
rect -564 215 -498 231
rect -446 265 -380 281
rect -446 231 -430 265
rect -396 231 -380 265
rect -446 215 -380 231
rect -328 265 -262 281
rect -328 231 -312 265
rect -278 231 -262 265
rect -328 215 -262 231
rect -210 265 -144 281
rect -210 231 -194 265
rect -160 231 -144 265
rect -210 215 -144 231
rect -92 265 -26 281
rect -92 231 -76 265
rect -42 231 -26 265
rect -92 215 -26 231
rect 26 265 92 281
rect 26 231 42 265
rect 76 231 92 265
rect 26 215 92 231
rect 144 265 210 281
rect 144 231 160 265
rect 194 231 210 265
rect 144 215 210 231
rect 262 265 328 281
rect 262 231 278 265
rect 312 231 328 265
rect 262 215 328 231
rect 380 265 446 281
rect 380 231 396 265
rect 430 231 446 265
rect 380 215 446 231
rect 498 265 564 281
rect 498 231 514 265
rect 548 231 564 265
rect 498 215 564 231
rect 616 265 682 281
rect 616 231 632 265
rect 666 231 682 265
rect 616 215 682 231
rect -679 193 -619 215
rect -561 193 -501 215
rect -443 193 -383 215
rect -325 193 -265 215
rect -207 193 -147 215
rect -89 193 -29 215
rect 29 193 89 215
rect 147 193 207 215
rect 265 193 325 215
rect 383 193 443 215
rect 501 193 561 215
rect 619 193 679 215
rect -679 87 -619 109
rect -561 87 -501 109
rect -443 87 -383 109
rect -325 87 -265 109
rect -207 87 -147 109
rect -89 87 -29 109
rect 29 87 89 109
rect 147 87 207 109
rect 265 87 325 109
rect 383 87 443 109
rect 501 87 561 109
rect 619 87 679 109
rect -682 71 -616 87
rect -682 37 -666 71
rect -632 37 -616 71
rect -682 21 -616 37
rect -564 71 -498 87
rect -564 37 -548 71
rect -514 37 -498 71
rect -564 21 -498 37
rect -446 71 -380 87
rect -446 37 -430 71
rect -396 37 -380 71
rect -446 21 -380 37
rect -328 71 -262 87
rect -328 37 -312 71
rect -278 37 -262 71
rect -328 21 -262 37
rect -210 71 -144 87
rect -210 37 -194 71
rect -160 37 -144 71
rect -210 21 -144 37
rect -92 71 -26 87
rect -92 37 -76 71
rect -42 37 -26 71
rect -92 21 -26 37
rect 26 71 92 87
rect 26 37 42 71
rect 76 37 92 71
rect 26 21 92 37
rect 144 71 210 87
rect 144 37 160 71
rect 194 37 210 71
rect 144 21 210 37
rect 262 71 328 87
rect 262 37 278 71
rect 312 37 328 71
rect 262 21 328 37
rect 380 71 446 87
rect 380 37 396 71
rect 430 37 446 71
rect 380 21 446 37
rect 498 71 564 87
rect 498 37 514 71
rect 548 37 564 71
rect 498 21 564 37
rect 616 71 682 87
rect 616 37 632 71
rect 666 37 682 71
rect 616 21 682 37
rect -682 -37 -616 -21
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -682 -87 -616 -71
rect -564 -37 -498 -21
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -564 -87 -498 -71
rect -446 -37 -380 -21
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -446 -87 -380 -71
rect -328 -37 -262 -21
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -328 -87 -262 -71
rect -210 -37 -144 -21
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -210 -87 -144 -71
rect -92 -37 -26 -21
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect -92 -87 -26 -71
rect 26 -37 92 -21
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 26 -87 92 -71
rect 144 -37 210 -21
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 144 -87 210 -71
rect 262 -37 328 -21
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 262 -87 328 -71
rect 380 -37 446 -21
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 380 -87 446 -71
rect 498 -37 564 -21
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 498 -87 564 -71
rect 616 -37 682 -21
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 616 -87 682 -71
rect -679 -109 -619 -87
rect -561 -109 -501 -87
rect -443 -109 -383 -87
rect -325 -109 -265 -87
rect -207 -109 -147 -87
rect -89 -109 -29 -87
rect 29 -109 89 -87
rect 147 -109 207 -87
rect 265 -109 325 -87
rect 383 -109 443 -87
rect 501 -109 561 -87
rect 619 -109 679 -87
rect -679 -215 -619 -193
rect -561 -215 -501 -193
rect -443 -215 -383 -193
rect -325 -215 -265 -193
rect -207 -215 -147 -193
rect -89 -215 -29 -193
rect 29 -215 89 -193
rect 147 -215 207 -193
rect 265 -215 325 -193
rect 383 -215 443 -193
rect 501 -215 561 -193
rect 619 -215 679 -193
rect -682 -231 -616 -215
rect -682 -265 -666 -231
rect -632 -265 -616 -231
rect -682 -281 -616 -265
rect -564 -231 -498 -215
rect -564 -265 -548 -231
rect -514 -265 -498 -231
rect -564 -281 -498 -265
rect -446 -231 -380 -215
rect -446 -265 -430 -231
rect -396 -265 -380 -231
rect -446 -281 -380 -265
rect -328 -231 -262 -215
rect -328 -265 -312 -231
rect -278 -265 -262 -231
rect -328 -281 -262 -265
rect -210 -231 -144 -215
rect -210 -265 -194 -231
rect -160 -265 -144 -231
rect -210 -281 -144 -265
rect -92 -231 -26 -215
rect -92 -265 -76 -231
rect -42 -265 -26 -231
rect -92 -281 -26 -265
rect 26 -231 92 -215
rect 26 -265 42 -231
rect 76 -265 92 -231
rect 26 -281 92 -265
rect 144 -231 210 -215
rect 144 -265 160 -231
rect 194 -265 210 -231
rect 144 -281 210 -265
rect 262 -231 328 -215
rect 262 -265 278 -231
rect 312 -265 328 -231
rect 262 -281 328 -265
rect 380 -231 446 -215
rect 380 -265 396 -231
rect 430 -265 446 -231
rect 380 -281 446 -265
rect 498 -231 564 -215
rect 498 -265 514 -231
rect 548 -265 564 -231
rect 498 -281 564 -265
rect 616 -231 682 -215
rect 616 -265 632 -231
rect 666 -265 682 -231
rect 616 -281 682 -265
<< polycont >>
rect -666 231 -632 265
rect -548 231 -514 265
rect -430 231 -396 265
rect -312 231 -278 265
rect -194 231 -160 265
rect -76 231 -42 265
rect 42 231 76 265
rect 160 231 194 265
rect 278 231 312 265
rect 396 231 430 265
rect 514 231 548 265
rect 632 231 666 265
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect -666 -265 -632 -231
rect -548 -265 -514 -231
rect -430 -265 -396 -231
rect -312 -265 -278 -231
rect -194 -265 -160 -231
rect -76 -265 -42 -231
rect 42 -265 76 -231
rect 160 -265 194 -231
rect 278 -265 312 -231
rect 396 -265 430 -231
rect 514 -265 548 -231
rect 632 -265 666 -231
<< locali >>
rect -839 333 -743 367
rect 743 333 839 367
rect -839 271 -805 333
rect 805 271 839 333
rect -682 231 -666 265
rect -632 231 -616 265
rect -564 231 -548 265
rect -514 231 -498 265
rect -446 231 -430 265
rect -396 231 -380 265
rect -328 231 -312 265
rect -278 231 -262 265
rect -210 231 -194 265
rect -160 231 -144 265
rect -92 231 -76 265
rect -42 231 -26 265
rect 26 231 42 265
rect 76 231 92 265
rect 144 231 160 265
rect 194 231 210 265
rect 262 231 278 265
rect 312 231 328 265
rect 380 231 396 265
rect 430 231 446 265
rect 498 231 514 265
rect 548 231 564 265
rect 616 231 632 265
rect 666 231 682 265
rect -725 181 -691 197
rect -725 105 -691 121
rect -607 181 -573 197
rect -607 105 -573 121
rect -489 181 -455 197
rect -489 105 -455 121
rect -371 181 -337 197
rect -371 105 -337 121
rect -253 181 -219 197
rect -253 105 -219 121
rect -135 181 -101 197
rect -135 105 -101 121
rect -17 181 17 197
rect -17 105 17 121
rect 101 181 135 197
rect 101 105 135 121
rect 219 181 253 197
rect 219 105 253 121
rect 337 181 371 197
rect 337 105 371 121
rect 455 181 489 197
rect 455 105 489 121
rect 573 181 607 197
rect 573 105 607 121
rect 691 181 725 197
rect 691 105 725 121
rect -682 37 -666 71
rect -632 37 -616 71
rect -564 37 -548 71
rect -514 37 -498 71
rect -446 37 -430 71
rect -396 37 -380 71
rect -328 37 -312 71
rect -278 37 -262 71
rect -210 37 -194 71
rect -160 37 -144 71
rect -92 37 -76 71
rect -42 37 -26 71
rect 26 37 42 71
rect 76 37 92 71
rect 144 37 160 71
rect 194 37 210 71
rect 262 37 278 71
rect 312 37 328 71
rect 380 37 396 71
rect 430 37 446 71
rect 498 37 514 71
rect 548 37 564 71
rect 616 37 632 71
rect 666 37 682 71
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 616 -71 632 -37
rect 666 -71 682 -37
rect -725 -121 -691 -105
rect -725 -197 -691 -181
rect -607 -121 -573 -105
rect -607 -197 -573 -181
rect -489 -121 -455 -105
rect -489 -197 -455 -181
rect -371 -121 -337 -105
rect -371 -197 -337 -181
rect -253 -121 -219 -105
rect -253 -197 -219 -181
rect -135 -121 -101 -105
rect -135 -197 -101 -181
rect -17 -121 17 -105
rect -17 -197 17 -181
rect 101 -121 135 -105
rect 101 -197 135 -181
rect 219 -121 253 -105
rect 219 -197 253 -181
rect 337 -121 371 -105
rect 337 -197 371 -181
rect 455 -121 489 -105
rect 455 -197 489 -181
rect 573 -121 607 -105
rect 573 -197 607 -181
rect 691 -121 725 -105
rect 691 -197 725 -181
rect -682 -265 -666 -231
rect -632 -265 -616 -231
rect -564 -265 -548 -231
rect -514 -265 -498 -231
rect -446 -265 -430 -231
rect -396 -265 -380 -231
rect -328 -265 -312 -231
rect -278 -265 -262 -231
rect -210 -265 -194 -231
rect -160 -265 -144 -231
rect -92 -265 -76 -231
rect -42 -265 -26 -231
rect 26 -265 42 -231
rect 76 -265 92 -231
rect 144 -265 160 -231
rect 194 -265 210 -231
rect 262 -265 278 -231
rect 312 -265 328 -231
rect 380 -265 396 -231
rect 430 -265 446 -231
rect 498 -265 514 -231
rect 548 -265 564 -231
rect 616 -265 632 -231
rect 666 -265 682 -231
rect -839 -333 -805 -271
rect 805 -333 839 -271
rect -839 -367 -743 -333
rect 743 -367 839 -333
<< viali >>
rect -666 231 -632 265
rect -548 231 -514 265
rect -430 231 -396 265
rect -312 231 -278 265
rect -194 231 -160 265
rect -76 231 -42 265
rect 42 231 76 265
rect 160 231 194 265
rect 278 231 312 265
rect 396 231 430 265
rect 514 231 548 265
rect 632 231 666 265
rect -725 121 -691 181
rect -607 121 -573 181
rect -489 121 -455 181
rect -371 121 -337 181
rect -253 121 -219 181
rect -135 121 -101 181
rect -17 121 17 181
rect 101 121 135 181
rect 219 121 253 181
rect 337 121 371 181
rect 455 121 489 181
rect 573 121 607 181
rect 691 121 725 181
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect -725 -181 -691 -121
rect -607 -181 -573 -121
rect -489 -181 -455 -121
rect -371 -181 -337 -121
rect -253 -181 -219 -121
rect -135 -181 -101 -121
rect -17 -181 17 -121
rect 101 -181 135 -121
rect 219 -181 253 -121
rect 337 -181 371 -121
rect 455 -181 489 -121
rect 573 -181 607 -121
rect 691 -181 725 -121
rect -666 -265 -632 -231
rect -548 -265 -514 -231
rect -430 -265 -396 -231
rect -312 -265 -278 -231
rect -194 -265 -160 -231
rect -76 -265 -42 -231
rect 42 -265 76 -231
rect 160 -265 194 -231
rect 278 -265 312 -231
rect 396 -265 430 -231
rect 514 -265 548 -231
rect 632 -265 666 -231
<< metal1 >>
rect -678 265 -620 271
rect -678 231 -666 265
rect -632 231 -620 265
rect -678 225 -620 231
rect -560 265 -502 271
rect -560 231 -548 265
rect -514 231 -502 265
rect -560 225 -502 231
rect -442 265 -384 271
rect -442 231 -430 265
rect -396 231 -384 265
rect -442 225 -384 231
rect -324 265 -266 271
rect -324 231 -312 265
rect -278 231 -266 265
rect -324 225 -266 231
rect -206 265 -148 271
rect -206 231 -194 265
rect -160 231 -148 265
rect -206 225 -148 231
rect -88 265 -30 271
rect -88 231 -76 265
rect -42 231 -30 265
rect -88 225 -30 231
rect 30 265 88 271
rect 30 231 42 265
rect 76 231 88 265
rect 30 225 88 231
rect 148 265 206 271
rect 148 231 160 265
rect 194 231 206 265
rect 148 225 206 231
rect 266 265 324 271
rect 266 231 278 265
rect 312 231 324 265
rect 266 225 324 231
rect 384 265 442 271
rect 384 231 396 265
rect 430 231 442 265
rect 384 225 442 231
rect 502 265 560 271
rect 502 231 514 265
rect 548 231 560 265
rect 502 225 560 231
rect 620 265 678 271
rect 620 231 632 265
rect 666 231 678 265
rect 620 225 678 231
rect -731 181 -685 193
rect -731 121 -725 181
rect -691 121 -685 181
rect -731 109 -685 121
rect -613 181 -567 193
rect -613 121 -607 181
rect -573 121 -567 181
rect -613 109 -567 121
rect -495 181 -449 193
rect -495 121 -489 181
rect -455 121 -449 181
rect -495 109 -449 121
rect -377 181 -331 193
rect -377 121 -371 181
rect -337 121 -331 181
rect -377 109 -331 121
rect -259 181 -213 193
rect -259 121 -253 181
rect -219 121 -213 181
rect -259 109 -213 121
rect -141 181 -95 193
rect -141 121 -135 181
rect -101 121 -95 181
rect -141 109 -95 121
rect -23 181 23 193
rect -23 121 -17 181
rect 17 121 23 181
rect -23 109 23 121
rect 95 181 141 193
rect 95 121 101 181
rect 135 121 141 181
rect 95 109 141 121
rect 213 181 259 193
rect 213 121 219 181
rect 253 121 259 181
rect 213 109 259 121
rect 331 181 377 193
rect 331 121 337 181
rect 371 121 377 181
rect 331 109 377 121
rect 449 181 495 193
rect 449 121 455 181
rect 489 121 495 181
rect 449 109 495 121
rect 567 181 613 193
rect 567 121 573 181
rect 607 121 613 181
rect 567 109 613 121
rect 685 181 731 193
rect 685 121 691 181
rect 725 121 731 181
rect 685 109 731 121
rect -678 71 -620 77
rect -678 37 -666 71
rect -632 37 -620 71
rect -678 31 -620 37
rect -560 71 -502 77
rect -560 37 -548 71
rect -514 37 -502 71
rect -560 31 -502 37
rect -442 71 -384 77
rect -442 37 -430 71
rect -396 37 -384 71
rect -442 31 -384 37
rect -324 71 -266 77
rect -324 37 -312 71
rect -278 37 -266 71
rect -324 31 -266 37
rect -206 71 -148 77
rect -206 37 -194 71
rect -160 37 -148 71
rect -206 31 -148 37
rect -88 71 -30 77
rect -88 37 -76 71
rect -42 37 -30 71
rect -88 31 -30 37
rect 30 71 88 77
rect 30 37 42 71
rect 76 37 88 71
rect 30 31 88 37
rect 148 71 206 77
rect 148 37 160 71
rect 194 37 206 71
rect 148 31 206 37
rect 266 71 324 77
rect 266 37 278 71
rect 312 37 324 71
rect 266 31 324 37
rect 384 71 442 77
rect 384 37 396 71
rect 430 37 442 71
rect 384 31 442 37
rect 502 71 560 77
rect 502 37 514 71
rect 548 37 560 71
rect 502 31 560 37
rect 620 71 678 77
rect 620 37 632 71
rect 666 37 678 71
rect 620 31 678 37
rect -678 -37 -620 -31
rect -678 -71 -666 -37
rect -632 -71 -620 -37
rect -678 -77 -620 -71
rect -560 -37 -502 -31
rect -560 -71 -548 -37
rect -514 -71 -502 -37
rect -560 -77 -502 -71
rect -442 -37 -384 -31
rect -442 -71 -430 -37
rect -396 -71 -384 -37
rect -442 -77 -384 -71
rect -324 -37 -266 -31
rect -324 -71 -312 -37
rect -278 -71 -266 -37
rect -324 -77 -266 -71
rect -206 -37 -148 -31
rect -206 -71 -194 -37
rect -160 -71 -148 -37
rect -206 -77 -148 -71
rect -88 -37 -30 -31
rect -88 -71 -76 -37
rect -42 -71 -30 -37
rect -88 -77 -30 -71
rect 30 -37 88 -31
rect 30 -71 42 -37
rect 76 -71 88 -37
rect 30 -77 88 -71
rect 148 -37 206 -31
rect 148 -71 160 -37
rect 194 -71 206 -37
rect 148 -77 206 -71
rect 266 -37 324 -31
rect 266 -71 278 -37
rect 312 -71 324 -37
rect 266 -77 324 -71
rect 384 -37 442 -31
rect 384 -71 396 -37
rect 430 -71 442 -37
rect 384 -77 442 -71
rect 502 -37 560 -31
rect 502 -71 514 -37
rect 548 -71 560 -37
rect 502 -77 560 -71
rect 620 -37 678 -31
rect 620 -71 632 -37
rect 666 -71 678 -37
rect 620 -77 678 -71
rect -731 -121 -685 -109
rect -731 -181 -725 -121
rect -691 -181 -685 -121
rect -731 -193 -685 -181
rect -613 -121 -567 -109
rect -613 -181 -607 -121
rect -573 -181 -567 -121
rect -613 -193 -567 -181
rect -495 -121 -449 -109
rect -495 -181 -489 -121
rect -455 -181 -449 -121
rect -495 -193 -449 -181
rect -377 -121 -331 -109
rect -377 -181 -371 -121
rect -337 -181 -331 -121
rect -377 -193 -331 -181
rect -259 -121 -213 -109
rect -259 -181 -253 -121
rect -219 -181 -213 -121
rect -259 -193 -213 -181
rect -141 -121 -95 -109
rect -141 -181 -135 -121
rect -101 -181 -95 -121
rect -141 -193 -95 -181
rect -23 -121 23 -109
rect -23 -181 -17 -121
rect 17 -181 23 -121
rect -23 -193 23 -181
rect 95 -121 141 -109
rect 95 -181 101 -121
rect 135 -181 141 -121
rect 95 -193 141 -181
rect 213 -121 259 -109
rect 213 -181 219 -121
rect 253 -181 259 -121
rect 213 -193 259 -181
rect 331 -121 377 -109
rect 331 -181 337 -121
rect 371 -181 377 -121
rect 331 -193 377 -181
rect 449 -121 495 -109
rect 449 -181 455 -121
rect 489 -181 495 -121
rect 449 -193 495 -181
rect 567 -121 613 -109
rect 567 -181 573 -121
rect 607 -181 613 -121
rect 567 -193 613 -181
rect 685 -121 731 -109
rect 685 -181 691 -121
rect 725 -181 731 -121
rect 685 -193 731 -181
rect -678 -231 -620 -225
rect -678 -265 -666 -231
rect -632 -265 -620 -231
rect -678 -271 -620 -265
rect -560 -231 -502 -225
rect -560 -265 -548 -231
rect -514 -265 -502 -231
rect -560 -271 -502 -265
rect -442 -231 -384 -225
rect -442 -265 -430 -231
rect -396 -265 -384 -231
rect -442 -271 -384 -265
rect -324 -231 -266 -225
rect -324 -265 -312 -231
rect -278 -265 -266 -231
rect -324 -271 -266 -265
rect -206 -231 -148 -225
rect -206 -265 -194 -231
rect -160 -265 -148 -231
rect -206 -271 -148 -265
rect -88 -231 -30 -225
rect -88 -265 -76 -231
rect -42 -265 -30 -231
rect -88 -271 -30 -265
rect 30 -231 88 -225
rect 30 -265 42 -231
rect 76 -265 88 -231
rect 30 -271 88 -265
rect 148 -231 206 -225
rect 148 -265 160 -231
rect 194 -265 206 -231
rect 148 -271 206 -265
rect 266 -231 324 -225
rect 266 -265 278 -231
rect 312 -265 324 -231
rect 266 -271 324 -265
rect 384 -231 442 -225
rect 384 -265 396 -231
rect 430 -265 442 -231
rect 384 -271 442 -265
rect 502 -231 560 -225
rect 502 -265 514 -231
rect 548 -265 560 -231
rect 502 -271 560 -265
rect 620 -231 678 -225
rect 620 -265 632 -231
rect 666 -265 678 -231
rect 620 -271 678 -265
<< properties >>
string FIXED_BBOX -822 -350 822 350
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 0.420 l 0.3 m 2 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
