magic
tech sky130A
magscale 1 2
timestamp 1645633816
<< dnwell >>
rect -200 -400 3400 2600
<< nwell >>
rect -280 2394 3480 2680
rect -280 -194 6 2394
rect 3194 -194 3480 2394
rect -280 -480 3480 -194
<< nsubdiff >>
rect -243 2623 3443 2643
rect -243 2589 -163 2623
rect 3363 2589 3443 2623
rect -243 2569 3443 2589
rect -243 2563 -169 2569
rect -243 -363 -223 2563
rect -189 -363 -169 2563
rect -243 -369 -169 -363
rect 3369 2563 3443 2569
rect 3369 -363 3389 2563
rect 3423 -363 3443 2563
rect 3369 -369 3443 -363
rect -243 -389 3443 -369
rect -243 -423 -163 -389
rect 3363 -423 3443 -389
rect -243 -443 3443 -423
<< nsubdiffcont >>
rect -163 2589 3363 2623
rect -223 -363 -189 2563
rect 3389 -363 3423 2563
rect -163 -423 3363 -389
<< locali >>
rect -223 2589 -163 2623
rect 3363 2589 3423 2623
rect -223 2563 -189 2589
rect -223 -389 -189 -363
rect 3389 2563 3423 2589
rect 3389 -389 3423 -363
rect -223 -423 -163 -389
rect 3363 -423 3423 -389
<< metal1 >>
rect 320 2020 2880 2080
rect 400 1140 460 2020
rect 2720 1140 2780 2020
rect 320 1000 2880 1140
rect 400 120 460 1000
rect 2720 120 2780 1000
rect 320 60 2900 120
use sky130_fd_pr__nfet_01v8_lvt_ZZ3Y87  sky130_fd_pr__nfet_01v8_lvt_ZZ3Y87_0
timestamp 1645633816
transform 1 0 1604 0 1 1066
box -1457 -1119 1457 1119
<< end >>
