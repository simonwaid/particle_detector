magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< pwell >>
rect 1340 7260 1840 7380
rect 1300 6040 1800 6140
<< locali >>
rect -20 13340 12960 13420
rect -20 7380 60 13340
rect -20 7358 10260 7380
rect 12860 7358 12960 13340
rect -20 7260 12960 7358
rect -20 7240 1340 7260
rect 1820 7246 12960 7260
rect 1820 7240 10260 7246
rect -20 6160 60 7240
rect -20 6140 1340 6160
rect 1760 6154 10360 6160
rect 12860 6154 12960 7246
rect 1760 6140 12960 6154
rect -20 6040 12960 6140
rect -20 5320 60 6040
rect 10074 6030 12960 6040
rect -20 60 60 5100
rect 12860 5320 12960 6030
rect 12860 60 12960 5080
rect -20 -40 12960 60
<< viali >>
rect -20 5100 60 5320
rect 12860 5080 12960 5320
<< metal1 >>
rect 1380 7138 1470 7172
rect 2638 7138 2728 7172
rect 3896 7138 3986 7172
rect 5154 7138 5244 7172
rect 1370 6840 1380 7040
rect 1460 6840 1470 7040
rect 3890 6840 3900 7040
rect 3980 6840 3990 7040
rect 130 6460 140 6660
rect 200 6460 210 6660
rect 2650 6460 2660 6660
rect 2720 6460 2730 6660
rect 5150 6460 5160 6660
rect 5240 6460 5250 6660
rect 1380 6228 1470 6262
rect 2638 6228 2728 6262
rect 3896 6228 3986 6262
rect 5154 6228 5244 6262
rect -26 5320 66 5332
rect -30 5100 -20 5320
rect 60 5100 70 5320
rect -26 5088 66 5100
rect 5600 140 6000 13260
rect 11450 7138 11540 7172
rect 12708 7138 12952 7172
rect 6410 6840 6420 7040
rect 6500 6840 6510 7040
rect 10190 6860 10200 7060
rect 10280 6860 10290 7060
rect 12690 6880 12700 7080
rect 12780 6880 12790 7080
rect 11450 6340 11460 6540
rect 11540 6340 11550 6540
rect 12916 6262 12952 7138
rect 11450 6228 11540 6262
rect 12708 6228 12952 6262
rect 11444 5928 11534 5962
rect 12854 5320 12966 5332
rect 12850 5080 12860 5320
rect 12960 5080 13120 5320
rect 12854 5068 12966 5080
<< via1 >>
rect 1380 6840 1460 7040
rect 3900 6840 3980 7040
rect 140 6460 200 6660
rect 2660 6460 2720 6660
rect 5160 6460 5240 6660
rect -20 5100 60 5320
rect 6420 6840 6500 7040
rect 10200 6860 10280 7060
rect 12700 6880 12780 7080
rect 11460 6340 11540 6540
rect 12860 5080 12960 5320
<< metal2 >>
rect 11380 13120 11660 13130
rect 11380 13010 11660 13020
rect 11840 11900 12040 11910
rect 11840 11790 12040 11800
rect 11380 10680 11660 10690
rect 11380 10570 11660 10580
rect 11360 9460 11640 9470
rect 11360 9350 11640 9360
rect 1880 8960 2180 8970
rect 1880 8810 2180 8820
rect 12700 8740 13100 8940
rect 11840 8240 12040 8250
rect 11840 8130 12040 8140
rect 12700 7520 13220 7720
rect 10200 7080 12880 7100
rect 10200 7060 12700 7080
rect 1380 7040 1460 7050
rect 3900 7040 3980 7050
rect 6420 7040 6500 7050
rect 140 6840 1380 7040
rect 1460 7000 3900 7040
rect 1460 6880 1880 7000
rect 2180 6880 3900 7000
rect 1460 6840 3900 6880
rect 3980 6840 6420 7040
rect 6500 6840 6520 7040
rect 10280 7000 12700 7060
rect 10280 6900 11840 7000
rect 12040 6900 12700 7000
rect 10280 6880 12700 6900
rect 12780 6880 12880 7080
rect 10280 6860 12880 6880
rect 10200 6840 12880 6860
rect 1380 6830 1460 6840
rect 3900 6830 3980 6840
rect 6420 6830 6500 6840
rect 140 6660 200 6670
rect 2660 6660 2720 6670
rect 5160 6660 5240 6670
rect 200 6620 2660 6660
rect 200 6500 220 6620
rect 520 6500 2660 6620
rect 200 6460 2660 6500
rect 2720 6460 5160 6660
rect 5240 6460 6460 6660
rect 11340 6540 11660 6560
rect 11340 6500 11460 6540
rect 11540 6500 11660 6540
rect 140 6450 200 6460
rect 2660 6450 2720 6460
rect 5160 6450 5240 6460
rect 11340 6400 11360 6500
rect 11640 6400 11660 6500
rect 11340 6340 11460 6400
rect 11540 6340 11660 6400
rect 11460 6330 11540 6340
rect 12460 5840 12660 5850
rect 1460 5820 1720 5830
rect 12460 5710 12660 5720
rect 1460 5690 1720 5700
rect -20 5320 60 5330
rect 12860 5320 12960 5330
rect 60 5100 200 5320
rect 620 5280 920 5290
rect 11840 5260 12040 5270
rect 11840 5150 12040 5160
rect 620 5130 920 5140
rect 12700 5100 12860 5320
rect -20 5090 60 5100
rect 12860 5070 12960 5080
rect 1880 4640 2180 4650
rect 1880 4490 2180 4500
rect 11360 4000 11640 4010
rect 11360 3890 11640 3900
rect 11360 2800 11640 2810
rect 11360 2690 11640 2700
rect 11840 1580 12040 1590
rect 11840 1470 12040 1480
rect 11360 360 11640 370
rect 11360 250 11640 260
<< via2 >>
rect 11380 13020 11660 13120
rect 11840 11800 12040 11900
rect 11380 10580 11660 10680
rect 11360 9360 11640 9460
rect 1880 8820 2180 8960
rect 11840 8140 12040 8240
rect 1880 6880 2180 7000
rect 11840 6900 12040 7000
rect 220 6500 520 6620
rect 11360 6400 11460 6500
rect 11460 6400 11540 6500
rect 11540 6400 11640 6500
rect 1460 5700 1720 5820
rect 12460 5720 12660 5840
rect 620 5140 920 5280
rect 11840 5160 12040 5260
rect 1880 4500 2180 4640
rect 11360 3900 11640 4000
rect 11360 2700 11640 2800
rect 11840 1480 12040 1580
rect 11360 260 11640 360
<< metal3 >>
rect 11360 13125 11660 13140
rect 11360 13120 11670 13125
rect 11360 13020 11380 13120
rect 11660 13020 11670 13120
rect 11360 13015 11670 13020
rect 216 6625 526 9460
rect 210 6620 530 6625
rect 210 6500 220 6620
rect 520 6500 530 6620
rect 210 6495 530 6500
rect 216 3960 526 6495
rect 620 5285 920 11620
rect 11360 10685 11660 13015
rect 11830 11900 12050 11905
rect 11830 11800 11840 11900
rect 12040 11800 12050 11900
rect 11830 11795 12050 11800
rect 11360 10680 11670 10685
rect 11360 10580 11380 10680
rect 11660 10580 11670 10680
rect 11360 10575 11670 10580
rect 11360 9465 11660 10575
rect 11350 9460 11660 9465
rect 11350 9360 11360 9460
rect 11640 9360 11660 9460
rect 11350 9355 11660 9360
rect 1870 8960 2190 8965
rect 1870 8820 1880 8960
rect 2180 8820 2190 8960
rect 1870 8815 2190 8820
rect 1880 7005 2180 8815
rect 1870 7000 2190 7005
rect 1870 6880 1880 7000
rect 2180 6880 2190 7000
rect 1870 6875 2190 6880
rect 1440 5900 1720 6160
rect 1380 5825 1720 5900
rect 1380 5820 1730 5825
rect 1380 5700 1460 5820
rect 1720 5700 1730 5820
rect 1380 5695 1730 5700
rect 1380 5680 1720 5695
rect 1380 5660 1680 5680
rect 610 5280 930 5285
rect 610 5140 620 5280
rect 920 5140 930 5280
rect 610 5135 930 5140
rect 620 1560 920 5135
rect 1880 4645 2180 6875
rect 11360 6505 11660 9355
rect 11840 8245 12040 11795
rect 11830 8240 12050 8245
rect 11830 8140 11840 8240
rect 12040 8140 12050 8240
rect 11830 8135 12050 8140
rect 11840 7005 12040 8135
rect 11830 7000 12050 7005
rect 11830 6900 11840 7000
rect 12040 6900 12050 7000
rect 11830 6895 12050 6900
rect 11350 6500 11660 6505
rect 11350 6400 11360 6500
rect 11640 6400 11660 6500
rect 11350 6395 11660 6400
rect 1870 4640 2190 4645
rect 1870 4500 1880 4640
rect 2180 4500 2190 4640
rect 1870 4495 2190 4500
rect 11360 4005 11660 6395
rect 11840 5265 12040 6895
rect 11830 5260 12050 5265
rect 11830 5160 11840 5260
rect 12040 5160 12050 5260
rect 11830 5155 12050 5160
rect 11350 4000 11660 4005
rect 11350 3900 11360 4000
rect 11640 3900 11660 4000
rect 11350 3895 11660 3900
rect 11360 2805 11660 3895
rect 11350 2800 11660 2805
rect 11350 2700 11360 2800
rect 11640 2700 11660 2800
rect 11350 2695 11660 2700
rect 11360 365 11660 2695
rect 11840 1585 12040 5155
rect 12120 4500 12320 8880
rect 12460 5845 12660 8940
rect 12450 5840 12670 5845
rect 12450 5720 12460 5840
rect 12660 5720 12670 5840
rect 12450 5715 12670 5720
rect 12460 4940 12660 5715
rect 11830 1580 12050 1585
rect 11830 1480 11840 1580
rect 12040 1480 12050 1580
rect 11830 1475 12050 1480
rect 11350 360 11660 365
rect 11350 260 11360 360
rect 11640 260 11660 360
rect 11350 255 11650 260
use isource_ref_5transistors  isource_ref_5transistors_0
timestamp 1654760956
transform 1 0 0 0 1 0
box 0 0 12914 4940
use isource_ref_5transistors  isource_ref_5transistors_1
timestamp 1654760956
transform 1 0 0 0 -1 13400
box 0 0 12914 4940
use isource_ref_transistor  isource_ref_transistor_0
timestamp 1654760956
transform 1 0 493 0 1 4997
box -493 -117 12421 1103
use sky130_fd_pr__nfet_01v8_TV3VM6  sky130_fd_pr__nfet_01v8_TV3VM6_0
timestamp 1654760956
transform 1 0 3312 0 1 6700
box -3312 -610 3312 610
use sky130_fd_pr__nfet_01v8_WY4VMC  sky130_fd_pr__nfet_01v8_WY4VMC_0
timestamp 1654760956
transform 1 0 11495 0 1 6700
box -1425 -610 1425 610
<< end >>
