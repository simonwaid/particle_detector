* SPICE3 file created from tia_core.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_CDW43Z a_100_n50# a_n100_n138# a_n260_n224# a_n158_n50#
X0 a_100_n50# a_n100_n138# a_n158_n50# a_n260_n224# sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_F8VELN a_n513_n200# a_n129_n200# a_399_n288# a_63_n200#
+ a_n225_n200# a_495_222# a_111_222# a_n321_n200# a_207_n288# a_n33_n200# a_n369_n288#
+ a_n707_n374# a_303_222# a_n605_n200# a_447_n200# a_15_n288# a_n81_222# a_n177_n288#
+ a_n561_n288# a_543_n200# a_159_n200# a_n273_222# a_255_n200# a_351_n200# a_n417_n200#
+ a_n465_222#
X0 a_n33_n200# a_n81_222# a_n129_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_351_n200# a_303_222# a_255_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_255_n200# a_207_n288# a_159_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n321_n200# a_n369_n288# a_n417_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_543_n200# a_495_222# a_447_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_159_n200# a_111_222# a_63_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_n225_n200# a_n273_222# a_n321_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X7 a_447_n200# a_399_n288# a_351_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 a_n513_n200# a_n561_n288# a_n605_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X9 a_63_n200# a_15_n288# a_n33_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 a_n129_n200# a_n177_n288# a_n225_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 a_n417_n200# a_n465_222# a_n513_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_854667 a_n287_n200# a_745_n200# a_n487_n288# a_545_n288#
+ a_229_n200# a_n545_n200# a_29_n288# a_n745_n288# a_487_n200# a_n29_n200# a_n229_n288#
+ a_n905_n374# a_287_n288# a_n803_n200#
X0 a_745_n200# a_545_n288# a_487_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X1 a_487_n200# a_287_n288# a_229_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X2 a_n29_n200# a_n229_n288# a_n287_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X3 a_229_n200# a_29_n288# a_n29_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4 a_n545_n200# a_n745_n288# a_n803_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X5 a_n287_n200# a_n487_n288# a_n545_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
.ends

.subckt tia_cur_mirror m1_71_n690# a_122_42# m1_71_130# m1_167_370# VSUBS
Xsky130_fd_pr__nfet_01v8_F8VELN_0 m1_167_370# m1_167_370# a_122_42# m1_167_370# m1_71_130#
+ a_122_42# a_122_42# m1_167_370# a_122_42# m1_71_130# a_122_42# VSUBS a_122_42# m1_71_130#
+ m1_167_370# a_122_42# a_122_42# a_122_42# a_122_42# m1_71_130# m1_71_130# a_122_42#
+ m1_167_370# m1_71_130# m1_71_130# a_122_42# sky130_fd_pr__nfet_01v8_F8VELN
Xsky130_fd_pr__nfet_01v8_854667_0 m1_71_n690# m1_71_n690# a_122_42# a_122_42# m1_71_n690#
+ m1_71_130# a_122_42# a_122_42# m1_71_130# m1_71_130# a_122_42# VSUBS a_122_42# m1_71_n690#
+ sky130_fd_pr__nfet_01v8_854667
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ZRA4RB a_n523_21# a_n817_n597# a_n1156_n509# a_n523_n87#
+ a_n1209_531# a_608_n509# a_216_109# a_n862_n509# a_n621_n597# a_n1209_n597# a_n568_109#
+ a_n78_n509# a_706_109# a_653_21# a_412_n509# a_653_n87# a_n817_531# a_n327_21# a_n131_n87#
+ a_n78_109# a_n1254_n509# a_n1058_109# a_n1013_n597# a_706_n509# a_n176_109# a_359_n597#
+ a_314_109# a_n176_n509# a_947_531# a_261_n87# a_n960_n509# a_n425_531# a_1143_n597#
+ a_457_21# a_n1111_n87# a_510_n509# a_n666_109# a_804_109# a_65_21# a_163_n597# a_n229_n597#
+ a_n1356_n683# a_n1156_109# a_555_531# a_804_n509# a_n274_n509# a_n915_21# a_n274_109#
+ a_412_109# a_1098_n509# a_n719_n87# a_n33_n597# a_1098_109# a_163_531# a_n764_109#
+ a_902_109# a_n568_n509# a_n33_531# a_n131_21# a_n1013_531# a_118_n509# a_902_n509#
+ a_n1254_109# a_849_n87# a_n719_21# a_n327_n87# a_555_n597# a_n372_n509# a_n1111_21#
+ a_1196_n509# a_1143_531# a_n372_109# a_510_109# a_261_21# a_20_109# a_n621_531#
+ a_1196_109# a_n666_n509# a_1000_109# a_n425_n597# a_849_21# a_n862_109# a_457_n87#
+ a_216_n509# a_1000_n509# a_751_531# a_n470_n509# a_n1058_n509# a_118_109# a_n470_109#
+ a_n229_531# a_n915_n87# a_947_n597# a_n764_n509# a_20_n509# a_608_109# a_1045_21#
+ a_n960_109# a_314_n509# a_65_n87# a_359_531# a_751_n597# a_1045_n87#
X0 a_n274_109# a_n327_21# a_n372_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X1 a_n764_n509# a_n817_n597# a_n862_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X2 a_706_n509# a_653_n87# a_608_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X3 a_n568_109# a_n621_531# a_n666_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X4 a_n862_109# a_n915_21# a_n960_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X5 a_1196_n509# a_1143_n597# a_1098_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X6 a_1196_109# a_1143_531# a_1098_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X7 a_n1156_n509# a_n1209_n597# a_n1254_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X8 a_n960_109# a_n1013_531# a_n1058_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X9 a_412_109# a_359_531# a_314_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X10 a_n470_n509# a_n523_n87# a_n568_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X11 a_n372_n509# a_n425_n597# a_n470_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X12 a_314_n509# a_261_n87# a_216_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X13 a_706_109# a_653_21# a_608_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X14 a_n862_n509# a_n915_n87# a_n960_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X15 a_n78_109# a_n131_21# a_n176_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X16 a_1000_109# a_947_531# a_902_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X17 a_804_n509# a_751_n597# a_706_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X18 a_n372_109# a_n425_531# a_n470_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X19 a_118_n509# a_65_n87# a_20_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X20 a_n666_109# a_n719_21# a_n764_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X21 a_n78_n509# a_n131_n87# a_n176_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X22 a_n1058_109# a_n1111_21# a_n1156_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X23 a_n568_n509# a_n621_n597# a_n666_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X24 a_412_n509# a_359_n597# a_314_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X25 a_216_109# a_163_531# a_118_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X26 a_118_109# a_65_21# a_20_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X27 a_510_109# a_457_21# a_412_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X28 a_n960_n509# a_n1013_n597# a_n1058_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X29 a_902_n509# a_849_n87# a_804_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X30 a_804_109# a_751_531# a_706_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X31 a_n176_109# a_n229_531# a_n274_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X32 a_n176_n509# a_n229_n597# a_n274_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X33 a_n470_109# a_n523_21# a_n568_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X34 a_n764_109# a_n817_531# a_n862_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X35 a_n666_n509# a_n719_n87# a_n764_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X36 a_510_n509# a_457_n87# a_412_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X37 a_1098_109# a_1045_21# a_1000_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X38 a_608_n509# a_555_n597# a_510_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X39 a_20_109# a_n33_531# a_n78_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X40 a_n1156_109# a_n1209_531# a_n1254_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X41 a_1000_n509# a_947_n597# a_902_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X42 a_1098_n509# a_1045_n87# a_1000_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X43 a_314_109# a_261_21# a_216_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X44 a_n1058_n509# a_n1111_n87# a_n1156_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X45 a_608_109# a_555_531# a_510_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X46 a_n274_n509# a_n327_n87# a_n372_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X47 a_902_109# a_849_21# a_804_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X48 a_20_n509# a_n33_n597# a_n78_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X49 a_216_n509# a_163_n597# a_118_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
.ends

.subckt sky130_fd_pr__pfet_01v8_NZHYX4 a_n568_n518# a_n764_118# a_653_n615# a_n719_n615#
+ a_163_n87# a_n33_n87# a_118_n518# a_n372_n518# a_n523_n615# a_510_118# a_n372_118#
+ a_20_118# a_65_549# a_n666_n518# a_n621_n87# a_163_21# a_n523_549# a_216_n518# a_n470_n518#
+ w_n902_n737# a_118_118# a_n470_118# a_653_549# a_n131_549# a_20_n518# a_n764_n518#
+ a_n229_n87# a_n621_21# a_314_n518# a_608_118# a_65_n615# a_359_n87# a_n33_21# a_261_549#
+ a_608_n518# a_216_118# a_n425_21# a_412_n518# a_n78_n518# a_706_118# a_n568_118#
+ a_457_n615# a_n78_118# a_555_21# a_n719_549# a_706_n518# a_n229_21# a_314_118# a_n176_118#
+ a_n176_n518# a_261_n615# a_n327_n615# a_510_n518# a_n425_n87# a_n666_118# a_359_21#
+ a_n327_549# a_n131_n615# a_n274_n518# a_555_n87# a_457_549# a_412_118# a_n274_118#
X0 a_n666_n518# a_n719_n615# a_n764_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X1 a_510_n518# a_457_n615# a_412_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X2 a_20_118# a_n33_21# a_n78_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X3 a_608_n518# a_555_n87# a_510_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X4 a_314_118# a_261_549# a_216_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X5 a_608_118# a_555_21# a_510_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X6 a_n274_n518# a_n327_n615# a_n372_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X7 a_20_n518# a_n33_n87# a_n78_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X8 a_216_n518# a_163_n87# a_118_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X9 a_n274_118# a_n327_549# a_n372_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X10 a_706_n518# a_653_n615# a_608_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X11 a_n568_118# a_n621_21# a_n666_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X12 a_412_118# a_359_21# a_314_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X13 a_n470_n518# a_n523_n615# a_n568_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X14 a_n372_n518# a_n425_n87# a_n470_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15 a_314_n518# a_261_n615# a_216_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X16 a_706_118# a_653_549# a_608_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X17 a_n78_118# a_n131_549# a_n176_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X18 a_n372_118# a_n425_21# a_n470_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X19 a_118_n518# a_65_n615# a_20_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X20 a_n666_118# a_n719_549# a_n764_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X21 a_n78_n518# a_n131_n615# a_n176_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X22 a_n568_n518# a_n621_n87# a_n666_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X23 a_412_n518# a_359_n87# a_314_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X24 a_118_118# a_65_549# a_20_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X25 a_216_118# a_163_21# a_118_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X26 a_510_118# a_457_549# a_412_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X27 a_n176_118# a_n229_21# a_n274_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X28 a_n176_n518# a_n229_n87# a_n274_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X29 a_n470_118# a_n523_549# a_n568_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
.ends

.subckt rf_transistors m1_2957_359# m1_1943_755# m1_2041_n2774# m1_3839_995# m1_1257_995#
+ m1_1551_n2534# m1_2727_n2534# m1_3643_119# m1_1061_119# m1_1061_n1330# m1_865_995#
+ m1_2237_n1330# m1_571_n2534# m1_1453_n472# m1_1747_359# m1_2761_755# m1_1061_n1916#
+ m1_2237_n1916# m1_3021_n472# m1_767_n712# m1_669_119# m1_1943_n2156# m1_2139_n2534#
+ a_622_n800# m1_1649_n2774# m1_2565_359# m1_1551_755# m1_963_n2156# m1_3447_995#
+ m1_1943_n1090# m1_3251_119# m1_669_n2774# m1_963_n1090# m1_2825_n2774# m1_571_n712#
+ m1_669_n472# m1_1355_359# m1_1159_n712# m1_1845_n1330# m1_1355_n2156# m1_963_359#
+ m1_2041_119# m1_1943_n712# m1_2335_n712# m1_865_n1330# m1_1845_n1916# m1_2369_755#
+ m1_1355_n1090# m1_2531_n2156# m1_3741_755# m1_3055_995# m1_865_n1916# m1_1061_n2774#
+ m1_2237_n2774# m1_2531_n1090# m1_1747_n2534# m1_2859_119# m1_1845_995# m1_1257_n1330#
+ m1_3545_359# m1_1159_755# m1_767_n2534# m1_1845_n472# m1_2237_n472# m1_2923_n2534#
+ m1_767_755# m1_571_359# m1_1257_n1916# a_623_n2862# m1_2433_n1330# m1_1649_119#
+ m1_2663_995# a_622_n2244# m1_2433_n1916# m1_1159_n2534# m1_2467_119# m1_1453_995#
+ m1_2335_n2534# m1_2041_n472# m1_3349_755# a_623_658# m1_1845_n2774# m1_3153_359#
+ m1_963_n712# m1_1943_359# m1_865_n2774# m1_3839_119# m1_1257_119# m1_3021_n1330#
+ m1_865_119# m1_2727_n712# m1_1551_n2156# m1_2727_n2156# m1_2957_755# m1_2761_359#
+ m1_3021_n1916# m1_3643_995# m1_571_n2156# m1_1257_n2774# a_623_22# m1_1061_995#
+ m1_1551_n1090# m1_2727_n1090# m1_865_n472# m1_1355_n712# m1_2433_n2774# m1_1747_755#
+ m1_571_n1090# m1_1943_n2534# m1_1551_359# m1_2629_n472# m1_2531_n712# m1_3447_119#
+ m1_1453_n1330# m1_2629_n1330# m1_2139_n2156# m1_669_995# m1_963_n2534# w_623_22#
+ m1_1453_n1916# m1_2565_755# m1_2139_n1090# m1_2629_n1916# m1_1257_n472# m1_3251_995#
+ a_623_n908# a_2421_658# m1_2433_n472# m1_1355_n2534# m1_2369_359# m1_3741_359# m1_1355_755#
+ m1_3021_n2774# m1_3055_119# m1_963_755# m1_2041_995# m1_2531_n2534# a_2421_22# m1_2041_n1330#
+ m1_1845_119# m1_1061_n472# m1_1159_359# m1_1747_n2156# m1_767_359# m1_2041_n1916#
+ m1_2859_995# m1_767_n2156# m1_1747_n1090# m1_2923_n2156# m1_2663_119# m1_3545_755#
+ m1_1747_n712# m1_1453_n2774# m1_2139_n712# m1_767_n1090# m1_2629_n2774# m1_571_755#
+ m1_2923_n712# m1_2923_n1090# m1_1649_995# m1_1649_n1330# m1_1159_n2156# m1_1453_119#
+ m1_3349_359# m1_669_n1330# m1_1649_n1916# m1_1159_n1090# m1_2825_n1330# m1_2335_n2156#
+ m1_1551_n712# m1_1649_n472# m1_2467_995# m1_669_n1916# m1_3153_755# VSUBS m1_2825_n472#
+ m1_2335_n1090# m1_2825_n1916#
Xsky130_fd_pr__nfet_01v8_lvt_ZRA4RB_0 a_622_n2244# a_623_n2862# m1_669_n2774# a_623_n2862#
+ a_622_n2244# m1_2433_n2774# m1_2041_n1916# m1_963_n2534# a_623_n2862# a_623_n2862#
+ m1_1257_n1916# m1_1747_n2534# m1_2531_n2156# a_622_n2244# m1_2237_n2774# a_623_n2862#
+ a_622_n2244# a_622_n2244# a_623_n2862# m1_1747_n2156# m1_571_n2534# m1_767_n2156#
+ a_623_n2862# m1_2531_n2534# m1_1649_n1916# a_623_n2862# m1_2139_n2156# m1_1649_n2774#
+ a_622_n2244# a_623_n2862# m1_865_n2774# a_622_n2244# a_623_n2862# a_622_n2244# a_623_n2862#
+ m1_2335_n2534# m1_1159_n2156# m1_2629_n1916# a_622_n2244# a_623_n2862# a_623_n2862#
+ VSUBS m1_669_n1916# a_622_n2244# m1_2629_n2774# m1_1551_n2534# a_622_n2244# m1_1551_n2156#
+ m1_2237_n1916# m1_2923_n2534# a_623_n2862# a_623_n2862# m1_2923_n2156# a_622_n2244#
+ m1_1061_n1916# m1_2727_n2156# m1_1257_n2774# a_622_n2244# a_622_n2244# a_622_n2244#
+ m1_1943_n2534# m1_2727_n2534# m1_571_n2156# a_623_n2862# a_622_n2244# a_623_n2862#
+ a_623_n2862# m1_1453_n2774# a_622_n2244# m1_3021_n2774# a_622_n2244# m1_1453_n1916#
+ m1_2335_n2156# a_622_n2244# m1_1845_n1916# a_622_n2244# m1_3021_n1916# m1_1159_n2534#
+ m1_2825_n1916# a_623_n2862# a_622_n2244# m1_963_n2156# a_623_n2862# m1_2041_n2774#
+ m1_2825_n2774# a_622_n2244# m1_1355_n2534# m1_767_n2534# m1_1943_n2156# m1_1355_n2156#
+ a_622_n2244# a_623_n2862# a_623_n2862# m1_1061_n2774# m1_1845_n2774# m1_2433_n1916#
+ a_622_n2244# m1_865_n1916# m1_2139_n2534# a_623_n2862# a_622_n2244# a_623_n2862#
+ a_623_n2862# sky130_fd_pr__nfet_01v8_lvt_ZRA4RB
Xsky130_fd_pr__nfet_01v8_lvt_ZRA4RB_1 a_622_n800# a_623_n908# m1_669_n1330# a_623_n908#
+ a_622_n800# m1_2433_n1330# m1_2041_n472# m1_963_n1090# a_623_n908# a_623_n908# m1_1257_n472#
+ m1_1747_n1090# m1_2531_n712# a_622_n800# m1_2237_n1330# a_623_n908# a_622_n800#
+ a_622_n800# a_623_n908# m1_1747_n712# m1_571_n1090# m1_767_n712# a_623_n908# m1_2531_n1090#
+ m1_1649_n472# a_623_n908# m1_2139_n712# m1_1649_n1330# a_622_n800# a_623_n908# m1_865_n1330#
+ a_622_n800# a_623_n908# a_622_n800# a_623_n908# m1_2335_n1090# m1_1159_n712# m1_2629_n472#
+ a_622_n800# a_623_n908# a_623_n908# VSUBS m1_669_n472# a_622_n800# m1_2629_n1330#
+ m1_1551_n1090# a_622_n800# m1_1551_n712# m1_2237_n472# m1_2923_n1090# a_623_n908#
+ a_623_n908# m1_2923_n712# a_622_n800# m1_1061_n472# m1_2727_n712# m1_1257_n1330#
+ a_622_n800# a_622_n800# a_622_n800# m1_1943_n1090# m1_2727_n1090# m1_571_n712# a_623_n908#
+ a_622_n800# a_623_n908# a_623_n908# m1_1453_n1330# a_622_n800# m1_3021_n1330# a_622_n800#
+ m1_1453_n472# m1_2335_n712# a_622_n800# m1_1845_n472# a_622_n800# m1_3021_n472#
+ m1_1159_n1090# m1_2825_n472# a_623_n908# a_622_n800# m1_963_n712# a_623_n908# m1_2041_n1330#
+ m1_2825_n1330# a_622_n800# m1_1355_n1090# m1_767_n1090# m1_1943_n712# m1_1355_n712#
+ a_622_n800# a_623_n908# a_623_n908# m1_1061_n1330# m1_1845_n1330# m1_2433_n472#
+ a_622_n800# m1_865_n472# m1_2139_n1090# a_623_n908# a_622_n800# a_623_n908# a_623_n908#
+ sky130_fd_pr__nfet_01v8_lvt_ZRA4RB
Xsky130_fd_pr__pfet_01v8_NZHYX4_1 m1_767_359# m1_571_755# a_623_22# a_623_22# a_623_22#
+ a_623_22# m1_1453_119# m1_963_359# a_623_22# m1_1845_995# m1_963_755# m1_1355_755#
+ a_623_658# m1_669_119# a_623_22# a_623_658# a_623_658# m1_1551_359# m1_865_119#
+ w_623_22# m1_1453_995# m1_865_995# a_623_658# a_623_658# m1_1355_359# m1_571_359#
+ a_623_22# a_623_658# m1_1649_119# m1_1943_755# a_623_22# a_623_22# a_623_658# a_623_658#
+ m1_1943_359# m1_1551_755# a_623_658# m1_1747_359# m1_1257_119# m1_2041_995# m1_767_755#
+ a_623_22# m1_1257_995# a_623_658# a_623_658# m1_2041_119# a_623_658# m1_1649_995#
+ m1_1159_755# m1_1159_359# a_623_22# a_623_22# m1_1845_119# a_623_22# m1_669_995#
+ a_623_658# a_623_658# a_623_22# m1_1061_119# a_623_22# a_623_658# m1_1747_755# m1_1061_995#
+ sky130_fd_pr__pfet_01v8_NZHYX4
Xsky130_fd_pr__pfet_01v8_NZHYX4_2 m1_2565_359# m1_2369_755# a_2421_22# a_2421_22#
+ a_2421_22# a_2421_22# m1_3251_119# m1_2761_359# a_2421_22# m1_3643_995# m1_2761_755#
+ m1_3153_755# a_2421_658# m1_2467_119# a_2421_22# a_2421_658# a_2421_658# m1_3349_359#
+ m1_2663_119# w_623_22# m1_3251_995# m1_2663_995# a_2421_658# a_2421_658# m1_3153_359#
+ m1_2369_359# a_2421_22# a_2421_658# m1_3447_119# m1_3741_755# a_2421_22# a_2421_22#
+ a_2421_658# a_2421_658# m1_3741_359# m1_3349_755# a_2421_658# m1_3545_359# m1_3055_119#
+ m1_3839_995# m1_2565_755# a_2421_22# m1_3055_995# a_2421_658# a_2421_658# m1_3839_119#
+ a_2421_658# m1_3447_995# m1_2957_755# m1_2957_359# a_2421_22# a_2421_22# m1_3643_119#
+ a_2421_22# m1_2467_995# a_2421_658# a_2421_658# a_2421_22# m1_2859_119# a_2421_22#
+ a_2421_658# m1_3545_755# m1_2859_995# sky130_fd_pr__pfet_01v8_NZHYX4
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_ZWVPUJ m4_n2851_n1900# c2_n2751_n1800#
X0 c2_n2751_n1800# m4_n2851_n1900# sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_RRWALQ a_n1041_109# a_n1041_727# a_1119_1149# a_n1185_21#
+ a_n1229_109# a_n1229_727# a_n753_n509# a_879_n1127# a_n81_727# a_447_639# a_n369_n509#
+ a_687_n1127# a_975_n1127# a_n81_109# a_n129_531# a_351_n87# a_399_n1127# a_495_n1127#
+ a_783_n1127# a_n33_n87# a_399_727# a_303_n509# a_591_n1127# a_399_109# a_n513_n597#
+ a_n129_n597# a_n321_639# a_879_109# a_879_727# a_63_n597# a_n273_109# a_n273_727#
+ a_n1089_n597# a_735_21# a_447_531# a_n225_n87# a_n465_n509# a_n753_727# a_n753_109#
+ a_n225_1149# a_15_109# a_15_727# a_n705_n705# a_1167_n509# a_255_n705# a_n321_531#
+ a_927_1149# a_n1185_1149# a_591_109# a_591_727# a_15_n509# a_n609_21# a_1119_21#
+ a_639_639# a_543_n87# a_n561_n509# a_1071_109# a_1071_727# a_1119_n1215# a_n177_n509#
+ a_n993_21# a_n33_n1215# a_207_727# a_n897_639# a_n321_n597# a_111_n509# a_207_109#
+ a_879_n509# a_n513_639# a_n609_n1215# a_n417_n1215# a_n1229_n1127# a_n465_727# a_639_n597#
+ a_n1185_n1215# a_n465_109# a_1023_n597# a_n801_n1215# a_n225_n1215# a_639_531# a_n417_n87#
+ a_n1137_n509# a_n273_n509# a_351_21# a_n945_727# a_n945_109# a_n1331_n1301# a_n897_531#
+ a_975_n509# a_831_639# a_n513_531# a_n513_n705# a_n129_n705# a_735_1149# a_n33_1149#
+ a_783_727# a_927_n1215# a_783_109# a_735_n1215# a_159_n1215# a_735_n87# a_543_n1215#
+ a_n33_21# a_n225_21# a_63_n705# a_351_n1215# a_n1089_n705# a_927_21# a_n1089_639#
+ a_15_n1127# a_n993_n87# a_n177_727# a_n177_109# a_831_531# a_n705_639# a_687_n509#
+ a_n897_n597# a_1071_n509# a_n657_727# a_831_n597# a_n657_109# a_447_n597# a_n993_n1215#
+ a_n609_n87# a_n1137_727# a_n1137_109# a_1023_639# a_n1089_531# a_495_727# a_n993_1149#
+ a_495_109# a_n1137_n1127# a_n705_531# a_111_727# a_n81_n509# a_783_n509# a_111_109#
+ a_n849_n509# a_399_n509# a_n321_n705# a_n1041_n1127# a_975_727# a_543_1149# a_63_639#
+ a_975_109# a_n609_1149# a_159_1149# a_927_n87# a_639_n705# a_n1041_n509# a_1023_n705#
+ a_1023_531# a_n1185_n87# a_543_21# a_n369_727# a_n369_109# a_159_21# a_n801_n87#
+ a_n945_n509# a_495_n509# a_207_n1127# a_n849_109# a_63_531# a_n849_727# a_255_639#
+ a_303_n1127# a_111_n1127# a_n705_n597# a_255_n597# a_1167_n1127# a_n801_21# a_159_n87#
+ a_n81_n1127# a_n417_21# a_1071_n1127# a_687_727# a_n1229_n509# a_687_109# a_303_727#
+ a_n849_n1127# a_303_109# a_1167_727# a_591_n509# a_1167_109# a_n657_n509# a_n945_n1127#
+ a_n657_n1127# a_n369_n1127# a_n897_n705# a_255_531# a_n129_639# a_n801_1149# a_1119_n87#
+ a_n753_n1127# a_n465_n1127# a_n177_n1127# a_351_1149# a_n561_n1127# a_n561_727#
+ a_n417_1149# a_n273_n1127# a_n561_109# a_831_n705# a_207_n509# a_447_n705#
X0 a_111_727# a_63_639# a_15_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_15_109# a_n33_21# a_n81_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_1071_n509# a_1023_n597# a_975_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n81_727# a_n129_639# a_n177_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n273_727# a_n321_639# a_n369_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_n177_727# a_n225_1149# a_n273_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 a_399_n509# a_351_n87# a_303_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_399_n1127# a_351_n1215# a_303_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X8 a_111_109# a_63_531# a_15_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X9 a_n465_n509# a_n513_n597# a_n561_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_n81_109# a_n129_531# a_n177_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X11 a_879_n1127# a_831_n705# a_783_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_n273_109# a_n321_531# a_n369_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X13 a_687_n509# a_639_n597# a_591_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X14 a_1071_n1127# a_1023_n705# a_975_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X15 a_n177_109# a_n225_21# a_n273_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 a_n81_n1127# a_n129_n705# a_n177_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17 a_n753_n509# a_n801_n87# a_n849_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X18 a_495_n1127# a_447_n705# a_399_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X19 a_n657_n1127# a_n705_n705# a_n753_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X20 a_975_n509# a_927_n87# a_879_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X21 a_975_n1127# a_927_n1215# a_879_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 a_n1137_n1127# a_n1185_n1215# a_n1229_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X23 a_n81_n509# a_n129_n597# a_n177_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X24 a_15_n509# a_n33_n87# a_n81_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X25 a_591_n1127# a_543_n1215# a_495_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X26 a_n753_n1127# a_n801_n1215# a_n849_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X27 a_n369_n509# a_n417_n87# a_n465_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X28 a_n1041_n509# a_n1089_n597# a_n1137_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X29 a_15_n1127# a_n33_n1215# a_n81_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X30 a_n657_n509# a_n705_n597# a_n753_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X31 a_879_n509# a_831_n597# a_783_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X32 a_n945_n509# a_n993_n87# a_n1041_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X33 a_1167_n509# a_1119_n87# a_1071_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X34 a_1167_n1127# a_1119_n1215# a_1071_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X35 a_n177_n1127# a_n225_n1215# a_n273_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X36 a_303_n509# a_255_n597# a_207_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X37 a_n273_n509# a_n321_n597# a_n369_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X38 a_303_727# a_255_639# a_207_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X39 a_591_727# a_543_1149# a_495_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X40 a_591_n509# a_543_n87# a_495_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X41 a_783_727# a_735_1149# a_687_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X42 a_495_727# a_447_639# a_399_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X43 a_207_727# a_159_1149# a_111_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 a_207_n1127# a_159_n1215# a_111_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X45 a_111_n1127# a_63_n705# a_15_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 a_n273_n1127# a_n321_n705# a_n369_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X47 a_975_727# a_927_1149# a_879_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X48 a_687_727# a_639_639# a_591_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 a_399_727# a_351_1149# a_303_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 a_n369_n1127# a_n417_n1215# a_n465_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X51 a_879_727# a_831_639# a_783_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 a_687_n1127# a_639_n705# a_591_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X53 a_n1041_727# a_n1089_639# a_n1137_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X54 a_n849_n1127# a_n897_n705# a_n945_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X55 a_n1137_727# a_n1185_1149# a_n1229_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X56 a_n849_n509# a_n897_n597# a_n945_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X57 a_1071_727# a_1023_639# a_975_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X58 a_n561_727# a_n609_1149# a_n657_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X59 a_303_n1127# a_255_n705# a_207_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 a_1167_727# a_1119_1149# a_1071_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X61 a_n465_727# a_n513_639# a_n561_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X62 a_n753_727# a_n801_1149# a_n849_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X63 a_n945_727# a_n993_1149# a_n1041_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X64 a_207_n509# a_159_n87# a_111_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X65 a_591_109# a_543_21# a_495_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X66 a_303_109# a_255_531# a_207_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X67 a_n369_727# a_n417_1149# a_n465_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 a_n657_727# a_n705_639# a_n753_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X69 a_n465_n1127# a_n513_n705# a_n561_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X70 a_207_109# a_159_21# a_111_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 a_n849_727# a_n897_639# a_n945_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X72 a_783_n1127# a_735_n1215# a_687_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 a_n177_n509# a_n225_n87# a_n273_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 a_783_109# a_735_21# a_687_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X75 a_495_109# a_447_531# a_399_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X76 a_687_109# a_639_531# a_591_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X77 a_399_109# a_351_21# a_303_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 a_975_109# a_927_21# a_879_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X79 a_n945_n1127# a_n993_n1215# a_n1041_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X80 a_879_109# a_831_531# a_783_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 a_n1041_109# a_n1089_531# a_n1137_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X82 a_15_727# a_n33_1149# a_n81_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X83 a_495_n509# a_447_n597# a_399_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 a_n1137_109# a_n1185_21# a_n1229_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X85 a_n1137_n509# a_n1185_n87# a_n1229_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X86 a_1071_109# a_1023_531# a_975_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X87 a_n561_n1127# a_n609_n1215# a_n657_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 a_n1041_n1127# a_n1089_n705# a_n1137_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 a_n561_109# a_n609_21# a_n657_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X90 a_n561_n509# a_n609_n87# a_n657_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 a_1167_109# a_1119_21# a_1071_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X92 a_n465_109# a_n513_531# a_n561_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X93 a_n753_109# a_n801_21# a_n849_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X94 a_111_n509# a_63_n597# a_15_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 a_n369_109# a_n417_21# a_n465_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 a_n657_109# a_n705_531# a_n753_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 a_n945_109# a_n993_21# a_n1041_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X98 a_783_n509# a_735_n87# a_687_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X99 a_n849_109# a_n897_531# a_n945_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt dis_tran m1_1422_1633# m1_1038_1633# m1_174_1015# m1_2190_775# m1_1326_157#
+ m1_78_2011# m1_750_1393# m1_1806_775# m1_558_157# m1_366_1393# m1_462_2011# m1_2094_1015#
+ m1_1422_397# m1_270_1633# m1_1134_1015# m1_654_397# m1_2286_1393# m1_1710_1393#
+ m1_2382_2011# m1_1326_1393# m1_270_775# m1_1422_2011# m1_1038_775# m1_1038_2011#
+ m1_2190_1633# m1_942_2251# m1_750_157# m1_558_2251# m1_1230_1633# m1_1518_157# m1_1998_1633#
+ m1_2382_775# m1_174_1393# m1_1998_397# m1_2478_2251# m1_270_2011# m1_78_775# m1_1614_397#
+ m1_1902_2251# m1_1518_2251# m1_846_397# m1_90_1210# m1_1230_775# m1_2094_1393# m1_846_1633#
+ m1_1134_1393# m1_462_775# m1_2190_2011# m1_1710_157# m1_90_1830# m1_1230_2011# m1_2094_157#
+ m1_1998_2011# m1_942_157# m1_750_2251# m1_366_2251# m1_1806_1633# m1_942_1015# m1_2190_397#
+ m1_558_1015# m1_1806_397# m1_90_590# m1_2286_2251# m1_1710_2251# m1_1326_2251# m1_1422_775#
+ m1_174_157# m1_846_2011# m1_2478_1015# m1_90_2440# m1_654_775# m1_1902_1015# m1_1902_157#
+ m1_654_1633# m1_1518_1015# m1_2286_157# m1_270_397# m1_1038_397# m1_174_2251# m1_1806_2011#
+ m1_2382_397# m1_1614_1633# m1_750_1015# m1_366_1015# m1_1134_157# m1_2094_2251#
+ m1_942_1393# m1_1998_775# m1_558_1393# m1_78_1633# m1_1614_775# m1_78_397# m1_1134_2251#
+ m1_366_157# m1_654_2011# m1_2286_1015# m1_846_775# m1_90_70# m1_1710_1015# m1_1230_397#
+ m1_462_1633# m1_2478_157# m1_1326_1015# m1_2478_1393# m1_462_397# m1_1902_1393#
+ m1_1518_1393# m1_1614_2011# m1_2382_1633# VSUBS
Xsky130_fd_pr__nfet_01v8_RRWALQ_0 m1_270_1633# m1_270_2011# m1_90_2440# m1_90_1210#
+ m1_78_1633# m1_78_2011# m1_558_1015# m1_2190_397# m1_1230_2011# m1_90_1830# m1_942_1015#
+ m1_1998_397# m1_2286_157# m1_1230_1633# m1_90_1830# m1_90_1210# m1_1710_157# m1_1806_397#
+ m1_2094_157# m1_90_1210# m1_1710_2251# m1_1614_775# m1_1902_157# m1_1710_1393# m1_90_590#
+ m1_90_590# m1_90_1830# m1_2190_1633# m1_2190_2011# m1_90_590# m1_1038_1633# m1_1038_2011#
+ m1_90_590# m1_90_1210# m1_90_1830# m1_90_1210# m1_846_775# m1_558_2251# m1_558_1393#
+ m1_90_2440# m1_1326_1393# m1_1326_2251# m1_90_590# m1_2478_1015# m1_90_590# m1_90_1830#
+ m1_90_2440# m1_90_2440# m1_1902_1393# m1_1902_2251# m1_1326_1015# m1_90_1210# m1_90_1210#
+ m1_90_1830# m1_90_1210# m1_750_1015# m1_2382_1633# m1_2382_2011# m1_90_70# m1_1134_1015#
+ m1_90_1210# m1_90_70# m1_1518_2251# m1_90_1830# m1_90_590# m1_1422_775# m1_1518_1393#
+ m1_2190_775# m1_90_1830# m1_90_70# m1_90_70# m1_78_397# m1_846_2011# m1_90_590#
+ m1_90_70# m1_846_1633# m1_90_590# m1_90_70# m1_90_70# m1_90_1830# m1_90_1210# m1_174_1015#
+ m1_1038_775# m1_90_1210# m1_366_2251# m1_366_1393# VSUBS m1_90_1830# m1_2286_1015#
+ m1_90_1830# m1_90_1830# m1_90_590# m1_90_590# m1_90_2440# m1_90_2440# m1_2094_2251#
+ m1_90_70# m1_2094_1393# m1_90_70# m1_90_70# m1_90_1210# m1_90_70# m1_90_1210# m1_90_1210#
+ m1_90_590# m1_90_70# m1_90_590# m1_90_1210# m1_90_1830# m1_1326_157# m1_90_1210#
+ m1_1134_2251# m1_1134_1393# m1_90_1830# m1_90_1830# m1_1998_775# m1_90_590# m1_2382_775#
+ m1_654_2011# m1_90_590# m1_654_1633# m1_90_590# m1_90_70# m1_90_1210# m1_174_2251#
+ m1_174_1393# m1_90_1830# m1_90_1830# m1_1806_2011# m1_90_2440# m1_1806_1633# m1_174_157#
+ m1_90_1830# m1_1422_2011# m1_1230_775# m1_2094_1015# m1_1422_1633# m1_462_775# m1_1710_1015#
+ m1_90_590# m1_270_397# m1_2286_2251# m1_90_2440# m1_90_1830# m1_2286_1393# m1_90_2440#
+ m1_90_2440# m1_90_1210# m1_90_590# m1_270_775# m1_90_590# m1_90_1830# m1_90_1210#
+ m1_90_1210# m1_942_2251# m1_942_1393# m1_90_1210# m1_90_1210# m1_366_1015# m1_1806_775#
+ m1_1518_157# m1_462_1633# m1_90_1830# m1_462_2011# m1_90_1830# m1_1614_397# m1_1422_397#
+ m1_90_590# m1_90_590# m1_2478_157# m1_90_1210# m1_90_1210# m1_1230_397# m1_90_1210#
+ m1_2382_397# m1_1998_2011# m1_78_775# m1_1998_1633# m1_1614_2011# m1_462_397# m1_1614_1633#
+ m1_2478_2251# m1_1902_1015# m1_2478_1393# m1_654_775# m1_366_157# m1_654_397# m1_942_157#
+ m1_90_590# m1_90_1830# m1_90_1830# m1_90_2440# m1_90_1210# m1_558_157# m1_846_397#
+ m1_1134_157# m1_90_2440# m1_750_157# m1_750_2251# m1_90_2440# m1_1038_397# m1_750_1393#
+ m1_90_590# m1_1518_1015# m1_90_590# sky130_fd_pr__nfet_01v8_RRWALQ
.ends

.subckt sky130_fd_pr__pfet_01v8_GYVK57 a_n819_n200# a_n345_n200# a_29_n297# a_n129_n297#
+ a_187_n297# a_129_n200# a_n503_n200# a_n287_n297# a_345_n297# a_287_n200# a_n661_n200#
+ a_n445_n297# a_503_n297# a_445_n200# a_n603_n297# a_661_n297# w_n957_n419# a_603_n200#
+ a_n761_n297# a_761_n200# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_761_n200# a_661_n297# a_603_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2 a_287_n200# a_187_n297# a_129_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3 a_n345_n200# a_n445_n297# a_n503_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X4 a_129_n200# a_29_n297# a_n29_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X5 a_445_n200# a_345_n297# a_287_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X6 a_n503_n200# a_n603_n297# a_n661_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X7 a_n29_n200# a_n129_n297# a_n187_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8 a_603_n200# a_503_n297# a_445_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9 a_n661_n200# a_n761_n297# a_n819_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_62U3RB a_608_n509# a_216_109# a_163_n87# a_n33_n87#
+ a_n327_531# a_n866_n683# a_n78_n509# a_n568_109# a_412_n509# a_706_109# a_n78_109#
+ a_457_531# a_706_n509# a_65_n597# a_n621_n87# a_n176_n509# a_314_109# a_n176_109#
+ a_163_21# a_510_n509# a_n666_109# a_n229_n87# a_n621_21# a_n274_n509# a_457_n597#
+ a_412_109# a_n274_109# a_65_531# a_n523_531# a_359_n87# a_n33_21# a_n568_n509# a_261_n597#
+ a_n327_n597# a_n764_109# a_118_n509# a_n425_21# a_653_531# a_n131_531# a_n372_n509#
+ a_n131_n597# a_510_109# a_n372_109# a_20_109# a_555_21# a_n666_n509# a_261_531#
+ a_n229_21# a_216_n509# a_653_n597# a_n470_n509# a_n425_n87# a_n719_n597# a_118_109#
+ a_n470_109# a_359_21# a_20_n509# a_n764_n509# a_n523_n597# a_608_109# a_314_n509#
+ a_555_n87# a_n719_531#
X0 a_n274_109# a_n327_531# a_n372_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X1 a_706_n509# a_653_n597# a_608_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X2 a_n568_109# a_n621_21# a_n666_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X3 a_412_109# a_359_21# a_314_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X4 a_n470_n509# a_n523_n597# a_n568_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X5 a_n372_n509# a_n425_n87# a_n470_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X6 a_314_n509# a_261_n597# a_216_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X7 a_706_109# a_653_531# a_608_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X8 a_n78_109# a_n131_531# a_n176_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X9 a_n372_109# a_n425_21# a_n470_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X10 a_118_n509# a_65_n597# a_20_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X11 a_n666_109# a_n719_531# a_n764_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X12 a_n78_n509# a_n131_n597# a_n176_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X13 a_n568_n509# a_n621_n87# a_n666_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X14 a_412_n509# a_359_n87# a_314_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X15 a_216_109# a_163_21# a_118_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X16 a_118_109# a_65_531# a_20_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X17 a_510_109# a_457_531# a_412_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X18 a_n176_109# a_n229_21# a_n274_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X19 a_n176_n509# a_n229_n87# a_n274_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X20 a_n470_109# a_n523_531# a_n568_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X21 a_n666_n509# a_n719_n597# a_n764_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X22 a_510_n509# a_457_n597# a_412_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X23 a_608_n509# a_555_n87# a_510_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X24 a_20_109# a_n33_21# a_n78_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X25 a_314_109# a_261_531# a_216_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X26 a_608_109# a_555_21# a_510_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X27 a_n274_n509# a_n327_n597# a_n372_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X28 a_20_n509# a_n33_n87# a_n78_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X29 a_216_n509# a_163_n87# a_118_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
.ends

.subckt fb_transistor m1_6753_3028# m1_6285_4403# sky130_fd_pr__pfet_01v8_GYVK57_0/a_503_n297#
+ m1_6459_2410# m1_7145_3028# m1_5871_3268# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n761_n297#
+ m1_6263_3268# m1_7145_2650# m1_6753_2650# m1_6917_4403# m1_6263_2410# m1_5871_2410#
+ m1_7233_4403# w_5706_2166# sky130_fd_pr__pfet_01v8_GYVK57_0/a_661_n297# m1_6127_4163#
+ a_5923_2832# m1_6759_4163# m1_5969_3028# m1_7075_4163# sky130_fd_pr__pfet_01v8_GYVK57_0/a_29_n297#
+ m1_5969_2650# m1_6655_3268# m1_6601_4403# m1_7047_3268# m1_6165_3028# m1_7047_2410#
+ m1_6655_2410# m1_7341_3028# m1_6165_2650# m1_6443_4163# m1_7341_2650# m1_7391_4163#
+ sky130_fd_pr__pfet_01v8_GYVK57_0/a_n129_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n287_n297#
+ m1_5811_4163# m1_6557_3028# m1_6851_3268# m1_6067_3268# sky130_fd_pr__pfet_01v8_GYVK57_0/a_187_n297#
+ m1_6557_2650# m1_7243_3268# m1_6067_2410# m1_6361_3028# a_5923_3450# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n445_n297#
+ m1_7243_2410# m1_6851_2410# m1_6361_2650# sky130_fd_pr__pfet_01v8_GYVK57_0/a_345_n297#
+ m1_6949_3028# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n603_n297# m1_6949_2650# m1_6459_3268#
+ m1_5969_4403# dw_5500_1960#
Xsky130_fd_pr__pfet_01v8_GYVK57_0 m1_5811_4163# m1_6285_4403# sky130_fd_pr__pfet_01v8_GYVK57_0/a_29_n297#
+ sky130_fd_pr__pfet_01v8_GYVK57_0/a_n129_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_187_n297#
+ m1_6759_4163# m1_6127_4163# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n287_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_345_n297#
+ m1_6917_4403# m1_5969_4403# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n445_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_503_n297#
+ m1_7075_4163# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n603_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_661_n297#
+ dw_5500_1960# m1_7233_4403# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n761_n297# m1_7391_4163#
+ m1_6601_4403# m1_6443_4163# sky130_fd_pr__pfet_01v8_GYVK57
Xsky130_fd_pr__nfet_01v8_lvt_62U3RB_0 m1_7243_2410# m1_6851_3268# a_5923_2832# a_5923_2832#
+ a_5923_3450# w_5706_2166# m1_6557_2650# m1_6067_3268# m1_7047_2410# m1_7341_3028#
+ m1_6557_3028# a_5923_3450# m1_7341_2650# a_5923_2832# a_5923_2832# m1_6459_2410#
+ m1_6949_3028# m1_6459_3268# a_5923_3450# m1_7145_2650# m1_5969_3028# a_5923_2832#
+ a_5923_3450# m1_6361_2650# a_5923_2832# m1_7047_3268# m1_6361_3028# a_5923_3450#
+ a_5923_3450# a_5923_2832# a_5923_3450# m1_6067_2410# a_5923_2832# a_5923_2832# m1_5871_3268#
+ m1_6753_2650# a_5923_3450# a_5923_3450# a_5923_3450# m1_6263_2410# a_5923_2832#
+ m1_7145_3028# m1_6263_3268# m1_6655_3268# a_5923_3450# m1_5969_2650# a_5923_3450#
+ a_5923_3450# m1_6851_2410# a_5923_2832# m1_6165_2650# a_5923_2832# a_5923_2832#
+ m1_6753_3028# m1_6165_3028# a_5923_3450# m1_6655_2410# m1_5871_2410# a_5923_2832#
+ m1_7243_3268# m1_6949_2650# a_5923_2832# a_5923_3450# sky130_fd_pr__nfet_01v8_lvt_62U3RB
.ends

.subckt tia_one_tia m1_n1960_n3240# m1_1850_2290# m2_1800_2380# tia_cur_mirror_0/m1_71_130#
+ w_1686_386# w_1650_2620# tia_cur_mirror_0/a_122_42# m2_n1840_n2910# VSUBS m1_1540_1550#
Xtia_cur_mirror_0 VSUBS tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# w_1686_386#
+ VSUBS tia_cur_mirror
Xrf_transistors_0 m1_1540_1550# m1_1540_1550# m2_n1840_n2910# w_1650_2620# w_1650_2620#
+ m1_1540_1550# m1_1540_1550# w_1650_2620# w_1650_2620# m2_n1840_n2910# w_1650_2620#
+ m2_n1840_n2910# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m2_n1840_n2910#
+ m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550# w_1650_2620# m1_1540_1550# m1_1540_1550#
+ w_1686_386# m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m1_1540_1550# w_1650_2620#
+ m1_1540_1550# w_1650_2620# m2_n1840_n2910# m1_1540_1550# m2_n1840_n2910# m1_1540_1550#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# m1_1540_1550#
+ w_1650_2620# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550#
+ m1_1540_1550# m1_1540_1550# m1_1540_1550# w_1650_2620# m2_n1840_n2910# m2_n1840_n2910#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# w_1650_2620# w_1650_2620# m2_n1840_n2910#
+ m1_1540_1550# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550#
+ m1_1540_1550# m1_1540_1550# m2_n1840_n2910# w_1686_386# m2_n1840_n2910# w_1650_2620#
+ w_1650_2620# w_1686_386# m2_n1840_n2910# m1_1540_1550# w_1650_2620# w_1650_2620#
+ m1_1540_1550# m2_n1840_n2910# m1_1540_1550# w_1686_386# m2_n1840_n2910# m1_1540_1550#
+ m1_1540_1550# m1_1540_1550# m2_n1840_n2910# w_1650_2620# w_1650_2620# m2_n1840_n2910#
+ w_1650_2620# m1_1540_1550# m1_1540_1550# m1_1540_1550# m1_1540_1550# m1_1540_1550#
+ m2_n1840_n2910# w_1650_2620# m1_1540_1550# m2_n1840_n2910# w_1686_386# w_1650_2620#
+ m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# m2_n1840_n2910# m1_1540_1550#
+ m1_1540_1550# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# w_1650_2620#
+ m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550# w_1650_2620# m1_1540_1550# w_1650_2620#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m2_n1840_n2910# w_1650_2620#
+ w_1686_386# w_1686_386# m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m1_1540_1550#
+ m1_1540_1550# m2_n1840_n2910# w_1650_2620# m1_1540_1550# w_1650_2620# m1_1540_1550#
+ w_1686_386# m2_n1840_n2910# w_1650_2620# m2_n1840_n2910# m1_1540_1550# m1_1540_1550#
+ m1_1540_1550# m2_n1840_n2910# w_1650_2620# m1_1540_1550# m1_1540_1550# m1_1540_1550#
+ w_1650_2620# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# m1_1540_1550#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m1_1540_1550# w_1650_2620# m2_n1840_n2910#
+ m1_1540_1550# w_1650_2620# m1_1540_1550# m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# w_1650_2620# m2_n1840_n2910#
+ m1_1540_1550# VSUBS m2_n1840_n2910# m1_1540_1550# m2_n1840_n2910# rf_transistors
Xsky130_fd_pr__cap_mim_m3_2_ZWVPUJ_0 m2_n1840_n2910# w_1650_2620# sky130_fd_pr__cap_mim_m3_2_ZWVPUJ
Xdis_tran_0 m2_n1840_n2910# m2_n1840_n2910# VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910#
+ m2_n1840_n2910# m2_n1840_n2910# m2_n1840_n2910# VSUBS VSUBS VSUBS m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# m2_n1840_n2910# VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910#
+ m2_n1840_n2910# m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# m1_n1960_n3240# m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910# VSUBS m1_n1960_n3240#
+ m2_n1840_n2910# VSUBS m2_n1840_n2910# VSUBS VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910#
+ VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910#
+ m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910# m2_n1840_n2910# VSUBS VSUBS
+ VSUBS VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910# m2_n1840_n2910#
+ VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m1_n1960_n3240# VSUBS m2_n1840_n2910#
+ m2_n1840_n2910# VSUBS VSUBS VSUBS m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# m2_n1840_n2910#
+ VSUBS dis_tran
Xfb_transistor_0 w_1686_386# w_1650_2620# m1_1850_2290# m2_1800_2380# w_1686_386#
+ m2_1800_2380# m1_1850_2290# m2_1800_2380# w_1686_386# w_1686_386# w_1650_2620# m2_1800_2380#
+ m2_1800_2380# w_1650_2620# w_1686_386# m1_1850_2290# m2_1800_2380# m1_1540_1550#
+ m2_1800_2380# w_1686_386# m2_1800_2380# m1_1850_2290# w_1686_386# m2_1800_2380#
+ w_1650_2620# m2_1800_2380# w_1686_386# m2_1800_2380# m2_1800_2380# w_1686_386# w_1686_386#
+ m2_1800_2380# w_1686_386# m2_1800_2380# m1_1850_2290# m1_1850_2290# m2_1800_2380#
+ w_1686_386# m2_1800_2380# m2_1800_2380# m1_1850_2290# w_1686_386# m2_1800_2380#
+ m2_1800_2380# w_1686_386# m1_1540_1550# m1_1850_2290# m2_1800_2380# m2_1800_2380#
+ w_1686_386# m1_1850_2290# w_1686_386# m1_1850_2290# w_1686_386# m2_1800_2380# w_1650_2620#
+ w_1650_2620# fb_transistor
.ends

.subckt sky130_fd_pr__pfet_01v8_GCYTE7 a_100_n50# w_n296_n269# a_n158_n50# a_n100_n147#
X0 a_100_n50# a_n100_n147# a_n158_n50# w_n296_n269# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_J5CT7Z c1_n1550_n1200# m3_n1650_n1300#
X0 c1_n1550_n1200# m3_n1650_n1300# sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
.ends

.subckt sky130_fd_pr__cap_var_lvt_MZUN4J a_n2040_n588# w_1507_n618# w_n2173_n618#
+ w_n333_n618# a_n1120_n588# w_587_n618# w_n1253_n618# a_n200_n588# a_1640_n588# a_720_n588#
X0 a_n200_n588# w_n333_n618# w_n333_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X1 a_n1120_n588# w_n1253_n618# w_n1253_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X2 a_720_n588# w_587_n618# w_587_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X3 a_1640_n588# w_1507_n618# w_1507_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X4 a_n2040_n588# w_n2173_n618# w_n2173_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG#0 m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_SC2JGL a_15_n200# a_n177_n200# a_111_n200# a_159_n288#
+ a_63_222# a_n81_n200# a_n129_222# a_n269_n200# a_207_n200# a_n225_n288# a_n371_n374#
+ a_n33_n288#
X0 a_n81_n200# a_n129_222# a_n177_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_15_n200# a_n33_n288# a_n81_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X2 a_207_n200# a_159_n288# a_111_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n177_n200# a_n225_n288# a_n269_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X4 a_111_n200# a_63_222# a_15_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt tia_core VPP Out_2 Out_1 Disable_TIA Input I_Bias1 VN
Xsky130_fd_pr__nfet_01v8_CDW43Z_0 VN Disable_TIA VN Disable_TIA_B sky130_fd_pr__nfet_01v8_CDW43Z
Xtia_cur_mirror_0 VN I_Bias1 VM6D I_Bias1 VN tia_cur_mirror
Xtia_one_tia_0 Disable_TIA_B VN Out_2 VM5D Input VPP I_Bias1 VM28D VN Out_1 tia_one_tia
Xtia_one_tia_1 Disable_TIA_B VN VM31D VM36D VM39D VPP I_Bias1 VM40D VN Out_ref tia_one_tia
Xsky130_fd_pr__pfet_01v8_GCYTE7_0 VPP VPP Disable_TIA_B Disable_TIA sky130_fd_pr__pfet_01v8_GCYTE7
Xsky130_fd_pr__cap_mim_m3_1_J5CT7Z_1 VN I_Bias1 sky130_fd_pr__cap_mim_m3_1_J5CT7Z
Xsky130_fd_pr__cap_mim_m3_1_J5CT7Z_0 VN I_Bias1 sky130_fd_pr__cap_mim_m3_1_J5CT7Z
Xsky130_fd_pr__cap_var_lvt_MZUN4J_0 Disable_TIA_B VN VN VN Disable_TIA_B VN VN Disable_TIA_B
+ Disable_TIA_B Disable_TIA_B sky130_fd_pr__cap_var_lvt_MZUN4J
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_0 VN VPP sky130_fd_pr__cap_mim_m3_2_LJ5JLG#0
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_1 VN VPP sky130_fd_pr__cap_mim_m3_2_LJ5JLG#0
Xsky130_fd_pr__nfet_01v8_SC2JGL_0 VN VN I_Bias1 Disable_TIA Disable_TIA I_Bias1 Disable_TIA
+ I_Bias1 VN Disable_TIA VN Disable_TIA sky130_fd_pr__nfet_01v8_SC2JGL
.ends

