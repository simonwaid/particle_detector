* SPICE3 file created from isource.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_1_WXTTNJ#0 c1_n2050_n2000# m3_n2150_n2100#
X0 c1_n2050_n2000# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_834VMG a_2487_n400# a_n29_n400# a_n2487_n488# a_1229_n400#
+ a_n2647_n574# a_n2545_n400# a_n1229_n488# a_1287_n488# a_n1287_n400# a_29_n488#
X0 a_n29_n400# a_n1229_n488# a_n1287_n400# a_n2647_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X1 a_n1287_n400# a_n2487_n488# a_n2545_n400# a_n2647_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X2 a_1229_n400# a_29_n488# a_n29_n400# a_n2647_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
X3 a_2487_n400# a_1287_n488# a_1229_n400# a_n2647_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_26RGPZ a_n225_n909# a_n129_109# a_n369_21# a_n465_931#
+ a_447_109# a_399_21# a_n321_n909# a_n177_n87# a_n81_n997# a_n321_109# a_n509_109#
+ a_n33_n909# a_n509_n909# a_159_109# a_n369_n87# a_111_931# a_447_n909# a_351_109#
+ a_n33_109# a_n611_n1083# a_159_n909# a_303_n997# a_n225_109# a_303_931# a_n177_21#
+ a_255_n909# a_399_n87# a_n465_n997# a_207_21# a_351_n909# a_n417_n909# a_63_109#
+ a_n81_931# a_15_n87# a_15_21# a_111_n997# a_n417_109# a_n273_931# a_n129_n909# a_n273_n997#
+ a_255_109# a_207_n87# a_63_n909#
X0 a_351_n909# a_303_n997# a_255_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X1 a_n33_n909# a_n81_n997# a_n129_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X2 a_255_n909# a_207_n87# a_159_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X3 a_n33_109# a_n81_931# a_n129_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X4 a_n321_n909# a_n369_n87# a_n417_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X5 a_351_109# a_303_931# a_255_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X6 a_159_109# a_111_931# a_63_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X7 a_255_109# a_207_21# a_159_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8 a_447_109# a_399_21# a_351_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.24e+12p pd=8.62e+06u as=0p ps=0u w=4e+06u l=150000u
X9 a_n321_109# a_n369_21# a_n417_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X10 a_n417_109# a_n465_931# a_n509_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.24e+12p ps=8.62e+06u w=4e+06u l=150000u
X11 a_n225_109# a_n273_931# a_n321_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=0p ps=0u w=4e+06u l=150000u
X12 a_n129_109# a_n177_21# a_n225_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 a_159_n909# a_111_n997# a_63_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X14 a_n225_n909# a_n273_n997# a_n321_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=0p ps=0u w=4e+06u l=150000u
X15 a_447_n909# a_399_n87# a_351_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.24e+12p pd=8.62e+06u as=0p ps=0u w=4e+06u l=150000u
X16 a_63_n909# a_15_n87# a_n33_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X17 a_63_109# a_15_21# a_n33_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 a_n129_n909# a_n177_n87# a_n225_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 a_n417_n909# a_n465_n997# a_n509_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.24e+12p ps=8.62e+06u w=4e+06u l=150000u
.ends

.subckt isource_conv_tsmal m1_4500_6730# m1_4590_7330# m1_4410_6620# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_26RGPZ_0 m1_4590_7330# m1_4500_6730# m1_4410_6620# m1_4410_6620#
+ m1_4500_6730# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4410_6620# m1_4500_6730#
+ m1_4500_6730# m1_4590_7330# m1_4500_6730# m1_4590_7330# m1_4410_6620# m1_4410_6620#
+ m1_4500_6730# m1_4590_7330# m1_4590_7330# VSUBS m1_4590_7330# m1_4410_6620# m1_4590_7330#
+ m1_4410_6620# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4410_6620# m1_4410_6620#
+ m1_4590_7330# m1_4590_7330# m1_4500_6730# m1_4410_6620# m1_4410_6620# m1_4410_6620#
+ m1_4410_6620# m1_4590_7330# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4500_6730#
+ m1_4410_6620# m1_4500_6730# sky130_fd_pr__nfet_01v8_lvt_26RGPZ
.ends

.subckt sky130_fd_pr__nfet_01v8_HZ8P49 a_2487_n400# a_n6261_n488# a_n29_n400# a_5003_n400#
+ a_3803_n488# a_n2487_n488# a_n3803_n400# a_n6421_n574# a_1229_n400# a_n5003_n488#
+ a_2545_n488# a_n2545_n400# a_n1229_n488# a_5061_n488# a_n5061_n400# a_3745_n400#
+ a_1287_n488# a_6261_n400# a_n1287_n400# a_29_n488# a_n6319_n400# a_n3745_n488#
X0 a_6261_n400# a_5061_n488# a_5003_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X1 a_n29_n400# a_n1229_n488# a_n1287_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X2 a_n2545_n400# a_n3745_n488# a_n3803_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X3 a_n1287_n400# a_n2487_n488# a_n2545_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4 a_5003_n400# a_3803_n488# a_3745_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X5 a_n3803_n400# a_n5003_n488# a_n5061_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X6 a_1229_n400# a_29_n488# a_n29_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
X7 a_3745_n400# a_2545_n488# a_2487_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X8 a_n5061_n400# a_n6261_n488# a_n6319_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X9 a_2487_n400# a_1287_n488# a_1229_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
.ends

.subckt isource_ref_transistor m1_n370_110# m1_887_21# m1_890_680# VSUBS
Xsky130_fd_pr__nfet_01v8_HZ8P49_0 m1_890_680# m1_887_21# m1_890_680# m1_890_680# m1_887_21#
+ m1_887_21# m1_n370_110# VSUBS m1_n370_110# m1_887_21# m1_887_21# m1_890_680# m1_887_21#
+ m1_887_21# m1_890_680# m1_n370_110# m1_887_21# m1_n370_110# m1_n370_110# m1_887_21#
+ m1_n370_110# m1_887_21# sky130_fd_pr__nfet_01v8_HZ8P49
.ends

.subckt sky130_fd_pr__pfet_01v8_ACY9XJ#0#0 a_20_n918# a_20_118# a_n78_n918# a_n33_21#
+ a_n78_118# w_n216_n1137# a_n33_n1015#
X0 a_20_118# a_n33_21# a_n78_118# w_n216_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X1 a_20_n918# a_n33_n1015# a_n78_n918# w_n216_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
.ends

.subckt sky130_fd_pr__pfet_01v8_J24RLQ#0#0 a_n416_118# a_n100_n1015# a_358_118# a_n416_n918#
+ a_n674_118# a_n158_118# a_n100_21# a_158_n1015# a_n358_21# w_n812_n1137# a_158_21#
+ a_358_n918# a_416_n1015# a_n358_n1015# a_100_n918# a_n674_n918# a_n616_21# a_416_21#
+ a_n616_n1015# a_n158_n918# a_616_118# a_100_118# a_616_n918#
X0 a_100_118# a_n100_21# a_n158_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X1 a_616_n918# a_416_n1015# a_358_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X2 a_358_n918# a_158_n1015# a_100_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X3 a_616_118# a_416_21# a_358_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X4 a_100_n918# a_n100_n1015# a_n158_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X5 a_358_118# a_158_21# a_100_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 a_n416_118# a_n616_21# a_n674_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X7 a_n416_n918# a_n616_n1015# a_n674_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X8 a_n158_n918# a_n358_n1015# a_n416_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 a_n158_118# a_n358_21# a_n416_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
.ends

.subckt isource_cmirror#0 m1_0_1060# li_0_0# m1_110_820#
Xsky130_fd_pr__pfet_01v8_ACY9XJ_0 m1_250_820# m1_250_820# m1_110_820# m1_0_1060# m1_110_820#
+ li_0_0# m1_0_1060# sky130_fd_pr__pfet_01v8_ACY9XJ#0#0
Xsky130_fd_pr__pfet_01v8_J24RLQ_0 li_0_0# m1_0_1060# m1_250_820# li_0_0# m1_250_820#
+ m1_250_820# m1_0_1060# m1_0_1060# m1_0_1060# li_0_0# m1_0_1060# m1_250_820# m1_0_1060#
+ m1_0_1060# li_0_0# m1_250_820# m1_0_1060# m1_0_1060# m1_0_1060# m1_250_820# li_0_0#
+ li_0_0# li_0_0# sky130_fd_pr__pfet_01v8_J24RLQ#0#0
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_JAGHGM a_n1331_n1562# a_n671_1000# a_919_n1432#
+ a_389_n1432# a_n141_1000# a_919_1000# a_389_1000# a_n141_n1432# a_n1201_n1432# a_n1201_1000#
+ a_n671_n1432#
X0 a_n1201_n1432# a_n1201_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1 a_919_n1432# a_919_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X2 a_n671_n1432# a_n671_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3 a_n141_n1432# a_n141_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X4 a_389_n1432# a_389_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
.ends

.subckt isource_out m1_18730_12160# isource_cmirror_0/m1_0_1060# m1_21256_12488# m1_20970_12680#
+ li_23190_12600# VSUBS isource_conv_tsmal_0/m1_4500_6730#
Xsky130_fd_pr__nfet_01v8_834VMG_0 VSUBS VSUBS m1_21256_12488# m1_18730_12160# VSUBS
+ VSUBS m1_21256_12488# m1_21256_12488# m1_18730_12160# m1_21256_12488# sky130_fd_pr__nfet_01v8_834VMG
Xisource_conv_tsmal_0 isource_conv_tsmal_0/m1_4500_6730# m1_16760_11560# m1_20970_12680#
+ VSUBS isource_conv_tsmal
Xisource_ref_transistor_0 m1_18730_12160# m1_16760_11560# m1_20970_12680# VSUBS isource_ref_transistor
Xisource_cmirror_0 isource_cmirror_0/m1_0_1060# li_23190_12600# m1_20970_12680# isource_cmirror#0
Xisource_ref_transistor_1 m1_20970_12680# m1_16760_11560# m1_18730_12160# VSUBS isource_ref_transistor
Xsky130_fd_pr__res_xhigh_po_1p41_JAGHGM_0 VSUBS m1_23460_11560# VSUBS m1_24000_9140#
+ m1_23460_11560# m1_24520_11560# m1_24520_11560# m1_24000_9140# m1_22920_9140# m1_16760_11560#
+ m1_22920_9140# sky130_fd_pr__res_xhigh_po_1p41_JAGHGM
.ends

.subckt isource_conv_tsmal_nwell m1_4500_6730# m1_4590_7330# w_4356_6496# dw_4150_6290#
+ m1_4410_6620#
Xsky130_fd_pr__nfet_01v8_lvt_26RGPZ_0 m1_4590_7330# m1_4500_6730# m1_4410_6620# m1_4410_6620#
+ m1_4500_6730# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4410_6620# m1_4500_6730#
+ m1_4500_6730# m1_4590_7330# m1_4500_6730# m1_4590_7330# m1_4410_6620# m1_4410_6620#
+ m1_4500_6730# m1_4590_7330# m1_4590_7330# w_4356_6496# m1_4590_7330# m1_4410_6620#
+ m1_4590_7330# m1_4410_6620# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4410_6620#
+ m1_4410_6620# m1_4590_7330# m1_4590_7330# m1_4500_6730# m1_4410_6620# m1_4410_6620#
+ m1_4410_6620# m1_4410_6620# m1_4590_7330# m1_4410_6620# m1_4500_6730# m1_4410_6620#
+ m1_4500_6730# m1_4410_6620# m1_4500_6730# sky130_fd_pr__nfet_01v8_lvt_26RGPZ
.ends

.subckt sky130_fd_pr__pfet_01v8_QDYTZD a_n200_n147# a_n258_n50# w_n396_n269# a_200_n50#
X0 a_200_n50# a_n200_n147# a_n258_n50# w_n396_n269# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_U3V43Z a_n258_n50# a_n200_n138# a_n360_n224# a_200_n50#
X0 a_200_n50# a_n200_n138# a_n258_n50# a_n360_n224# sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_E9U3PA a_363_n400# a_114_n488# a_n29_n400# a_408_422#
+ a_n278_n488# a_461_n400# a_n127_n400# a_n180_422# a_n82_n488# a_16_422# a_n225_n400#
+ a_310_n488# a_n519_n400# a_69_n400# a_n323_n400# a_n474_n488# a_212_422# a_167_n400#
+ a_n376_422# a_n421_n400# a_265_n400# a_n621_n574#
X0 a_n421_n400# a_n474_n488# a_n519_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X1 a_461_n400# a_408_422# a_363_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X2 a_n127_n400# a_n180_422# a_n225_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X3 a_167_n400# a_114_n488# a_69_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X4 a_n225_n400# a_n278_n488# a_n323_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X5 a_265_n400# a_212_422# a_167_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=200000u
X6 a_69_n400# a_16_422# a_n29_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X7 a_n323_n400# a_n376_422# a_n421_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X8 a_n29_n400# a_n82_n488# a_n127_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X9 a_363_n400# a_310_n488# a_265_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
.ends

.subckt isource_startup li_2190_920# m1_360_100# sky130_fd_pr__nfet_01v8_U3V43Z_0/a_200_n50#
+ VSUBS
Xsky130_fd_pr__pfet_01v8_QDYTZD_1 m1_360_100# m1_330_800# li_2190_920# li_2190_920#
+ sky130_fd_pr__pfet_01v8_QDYTZD
Xsky130_fd_pr__nfet_01v8_U3V43Z_0 VSUBS m1_330_800# VSUBS sky130_fd_pr__nfet_01v8_U3V43Z_0/a_200_n50#
+ sky130_fd_pr__nfet_01v8_U3V43Z
Xsky130_fd_pr__nfet_01v8_lvt_E9U3PA_0 VSUBS m1_360_100# VSUBS m1_360_100# m1_360_100#
+ m1_330_800# m1_330_800# m1_360_100# m1_360_100# m1_360_100# VSUBS m1_360_100# m1_330_800#
+ m1_330_800# m1_330_800# m1_360_100# m1_360_100# VSUBS m1_360_100# VSUBS m1_330_800#
+ VSUBS sky130_fd_pr__nfet_01v8_lvt_E9U3PA
.ends

.subckt isource_ref_5transistors m2_12120_850# m1_12450_1060# m2_220_270# VSUBS
Xisource_ref_transistor_0 m2_220_270# m1_12450_1060# m2_12120_850# VSUBS isource_ref_transistor
Xisource_ref_transistor_1 VSUBS m1_12450_1060# m1_12450_1060# VSUBS isource_ref_transistor
Xisource_ref_transistor_3 m2_220_270# m1_12450_1060# m2_12120_850# VSUBS isource_ref_transistor
Xisource_ref_transistor_4 m2_220_270# m1_12450_1060# m2_12120_850# VSUBS isource_ref_transistor
.ends

.subckt sky130_fd_pr__nfet_01v8_TV3VM6 a_n658_n400# a_n3276_n574# a_n600_n488# a_n3174_n400#
+ a_1858_n400# a_n1858_n488# a_3116_n400# a_1916_n488# a_658_n488# a_600_n400# a_n1916_n400#
+ a_n3116_n488#
X0 a_1858_n400# a_658_n488# a_600_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X1 a_n658_n400# a_n1858_n488# a_n1916_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X2 a_n1916_n400# a_n3116_n488# a_n3174_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X3 a_3116_n400# a_1916_n488# a_1858_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
X4 a_600_n400# a_n600_n488# a_n658_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_WY4VMC a_n29_n400# a_1229_n400# a_n1229_n488# a_n1389_n574#
+ a_n1287_n400# a_29_n488#
X0 a_n29_n400# a_n1229_n488# a_n1287_n400# a_n1389_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X1 a_1229_n400# a_29_n488# a_n29_n400# a_n1389_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
.ends

.subckt isource_ref m2_12700_7520# m1_1370_6840# m1_12708_6228# m1_5600_140# m1_130_6460#
+ VSUBS
Xisource_ref_transistor_0 VSUBS m1_5600_140# m1_5600_140# VSUBS isource_ref_transistor
Xisource_ref_5transistors_0 m1_1370_6840# m1_5600_140# m1_130_6460# VSUBS isource_ref_5transistors
Xisource_ref_5transistors_1 m1_1370_6840# m1_5600_140# m1_130_6460# VSUBS isource_ref_5transistors
Xsky130_fd_pr__nfet_01v8_TV3VM6_0 m1_130_6460# VSUBS m1_5600_140# m1_130_6460# m1_130_6460#
+ m1_5600_140# m1_1370_6840# m1_5600_140# m1_5600_140# m1_1370_6840# m1_1370_6840#
+ m1_5600_140# sky130_fd_pr__nfet_01v8_TV3VM6
Xsky130_fd_pr__nfet_01v8_WY4VMC_0 m1_130_6460# VSUBS m1_12708_6228# VSUBS VSUBS m1_12708_6228#
+ sky130_fd_pr__nfet_01v8_WY4VMC
.ends

.subckt sky130_fd_pr__pfet_01v8_ACY9XJ#0 a_20_n918# a_20_118# a_n78_n918# a_n33_21#
+ a_n78_118# w_n216_n1137# a_n33_n1015#
X0 a_20_118# a_n33_21# a_n78_118# w_n216_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X1 a_20_n918# a_n33_n1015# a_n78_n918# w_n216_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
.ends

.subckt sky130_fd_pr__pfet_01v8_J24RLQ#0 a_n416_118# a_n100_n1015# a_358_118# a_n416_n918#
+ a_n674_118# a_n158_118# a_n100_21# a_158_n1015# a_n358_21# w_n812_n1137# a_158_21#
+ a_358_n918# a_416_n1015# a_n358_n1015# a_100_n918# a_n674_n918# a_n616_21# a_416_21#
+ a_n616_n1015# a_n158_n918# a_616_118# a_100_118# a_616_n918#
X0 a_100_118# a_n100_21# a_n158_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X1 a_616_n918# a_416_n1015# a_358_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X2 a_358_n918# a_158_n1015# a_100_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X3 a_616_118# a_416_21# a_358_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X4 a_100_n918# a_n100_n1015# a_n158_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X5 a_358_118# a_158_21# a_100_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 a_n416_118# a_n616_21# a_n674_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X7 a_n416_n918# a_n616_n1015# a_n674_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X8 a_n158_n918# a_n358_n1015# a_n416_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 a_n158_118# a_n358_21# a_n416_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
.ends

.subckt isource_cmirror m1_0_1060# li_0_0# m1_250_820# m1_110_820#
Xsky130_fd_pr__pfet_01v8_ACY9XJ_0 m1_250_820# m1_250_820# m1_110_820# m1_0_1060# m1_110_820#
+ li_0_0# m1_0_1060# sky130_fd_pr__pfet_01v8_ACY9XJ#0
Xsky130_fd_pr__pfet_01v8_J24RLQ_0 li_0_0# m1_0_1060# m1_250_820# li_0_0# m1_250_820#
+ m1_250_820# m1_0_1060# m1_0_1060# m1_0_1060# li_0_0# m1_0_1060# m1_250_820# m1_0_1060#
+ m1_0_1060# li_0_0# m1_250_820# m1_0_1060# m1_0_1060# m1_0_1060# m1_250_820# li_0_0#
+ li_0_0# li_0_0# sky130_fd_pr__pfet_01v8_J24RLQ#0
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_BQY2W7 a_n406_1000# a_n1996_1000# a_n1996_n1432#
+ a_654_n1432# a_1714_1000# a_1714_n1432# a_1184_n1432# a_n1466_1000# a_1184_1000#
+ a_n2126_n1562# a_n406_n1432# a_654_1000# a_n936_1000# a_n936_n1432# a_n1466_n1432#
+ a_124_n1432# a_124_1000#
X0 a_654_n1432# a_654_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1 a_124_n1432# a_124_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X2 a_n1996_n1432# a_n1996_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3 a_n1466_n1432# a_n1466_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X4 a_n936_n1432# a_n936_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X5 a_1714_n1432# a_1714_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X6 a_n406_n1432# a_n406_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X7 a_1184_n1432# a_1184_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_J2NVFM a_n406_1000# a_n406_n1432# a_124_n1432#
+ a_124_1000# a_n536_n1562#
X0 a_124_n1432# a_124_1000# a_n536_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1 a_n406_n1432# a_n406_1000# a_n536_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
.ends

.subckt isource_conv m1_4090_13100# m1_9600_7000# m1_4700_7820# m2_10060_7720# m1_5350_12620#
+ sky130_fd_pr__res_xhigh_po_1p41_BQY2W7_0/a_1714_n1432# li_9700_9140# VSUBS m1_4150_7820#
Xisource_cmirror_0 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_1 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_2 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_3 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_4 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_5 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xsky130_fd_pr__res_xhigh_po_1p41_BQY2W7_0 m1_6360_10260# m1_5300_10260# m1_4700_7820#
+ m1_7960_7820# m1_8480_10260# sky130_fd_pr__res_xhigh_po_1p41_BQY2W7_0/a_1714_n1432#
+ m1_7960_7820# m1_5300_10260# m1_8480_10260# VSUBS m1_6900_7820# m1_7420_10260# m1_6360_10260#
+ m1_5840_7820# m1_5840_7820# m1_6900_7820# m1_7420_10260# sky130_fd_pr__res_xhigh_po_1p41_BQY2W7
Xsky130_fd_pr__nfet_01v8_WY4VMC_2 m1_5350_12620# m1_4090_13100# m1_4150_7820# VSUBS
+ m1_4090_13100# m1_4150_7820# sky130_fd_pr__nfet_01v8_WY4VMC
Xsky130_fd_pr__res_xhigh_po_1p41_J2NVFM_0 m1_4160_10260# m1_4150_7820# m1_4700_7820#
+ m1_4160_10260# VSUBS sky130_fd_pr__res_xhigh_po_1p41_J2NVFM
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ZZ3Y87 a_n287_n909# a_n229_n997# a_n1003_n997#
+ a_229_109# a_n1061_n909# a_287_n997# a_n487_21# a_n1061_109# a_745_n909# a_n545_109#
+ a_287_21# a_n1261_21# a_1061_n997# a_487_109# a_n745_21# a_229_n909# a_n29_109#
+ a_1061_21# a_29_21# a_n487_n997# a_n1261_n997# a_545_21# a_n545_n909# a_n287_109#
+ a_545_n997# a_1003_n909# a_1003_109# a_n29_n909# a_803_21# a_487_n909# a_29_n997#
+ a_n229_21# a_n745_n997# a_n803_n909# a_n803_109# a_n1319_109# a_803_n997# a_1261_109#
+ a_n1003_21# a_n1421_n1083# a_1261_n909# a_745_109# a_n1319_n909#
X0 a_229_109# a_29_21# a_n29_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X1 a_1261_n909# a_1061_n997# a_1003_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X2 a_487_109# a_287_21# a_229_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=1e+06u
X3 a_n545_109# a_n745_21# a_n803_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X4 a_1261_109# a_1061_21# a_1003_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X5 a_n29_n909# a_n229_n997# a_n287_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X6 a_229_n909# a_29_n997# a_n29_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=1e+06u
X7 a_n1061_109# a_n1261_21# a_n1319_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X8 a_n287_109# a_n487_21# a_n545_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=1e+06u
X9 a_n545_n909# a_n745_n997# a_n803_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X10 a_n287_n909# a_n487_n997# a_n545_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11 a_n803_n909# a_n1003_n997# a_n1061_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X12 a_1003_109# a_803_21# a_745_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X13 a_n1061_n909# a_n1261_n997# a_n1319_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X14 a_1003_n909# a_803_n997# a_745_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X15 a_n803_109# a_n1003_21# a_n1061_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X16 a_745_n909# a_545_n997# a_487_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X17 a_n29_109# a_n229_21# a_n287_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X18 a_745_109# a_545_21# a_487_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X19 a_487_n909# a_287_n997# a_229_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
.ends

.subckt isource_diffamp dw_14640_n8120# w_14846_n7914# m1_15050_n7600# m1_14640_n6760#
+ m1_15310_n7040#
Xsky130_fd_pr__nfet_01v8_lvt_ZZ3Y87_0 m1_15050_n7600# m1_14640_n6760# m1_14640_n6760#
+ m1_15050_n7600# m1_15310_n7040# m1_14640_n6760# m1_14640_n6760# m1_15310_n7040#
+ m1_15050_n7600# m1_15310_n7040# m1_14640_n6760# m1_14640_n6760# m1_14640_n6760#
+ m1_15310_n7040# m1_14640_n6760# m1_15050_n7600# m1_15310_n7040# m1_14640_n6760#
+ m1_14640_n6760# m1_14640_n6760# m1_14640_n6760# m1_14640_n6760# m1_15310_n7040#
+ m1_15050_n7600# m1_14640_n6760# m1_15310_n7040# m1_15310_n7040# m1_15310_n7040#
+ m1_14640_n6760# m1_15310_n7040# m1_14640_n6760# m1_14640_n6760# m1_14640_n6760#
+ m1_15050_n7600# m1_15050_n7600# m1_15050_n7600# m1_14640_n6760# m1_15050_n7600#
+ m1_14640_n6760# w_14846_n7914# m1_15050_n7600# m1_15050_n7600# m1_15050_n7600# sky130_fd_pr__nfet_01v8_lvt_ZZ3Y87
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG#1 m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt isource VP I_ref VN
Xsky130_fd_pr__cap_mim_m3_1_WXTTNJ_0 VP VM8D sky130_fd_pr__cap_mim_m3_1_WXTTNJ#0
Xisource_out_0 VM3D VM8D VM3G VM22D VP VN I_ref isource_out
Xisource_conv_tsmal_nwell_0 VP VM12G VM12G VP VM14D isource_conv_tsmal_nwell
Xisource_startup_0 VP VM11D VM8D VN isource_startup
Xisource_ref_0 VM11D VM11D VM12G VM2D VM12D VN isource_ref
Xisource_cmirror_2 VM8D VP VM9D isource_cmirror#0
Xisource_cmirror_3 VM8D VP VM8D isource_cmirror#0
Xisource_conv_0 VN VM8D VM3G m2_19160_1520# VM14D VN VP VN VM12G isource_conv
Xisource_diffamp_0 VP VM11D VM11D VM9D VM8D isource_diffamp
Xisource_diffamp_1 VP VM2D VM2D VM9D VM9D isource_diffamp
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_0 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#1
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_1 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#1
.ends

