* SPICE3 file created from mpw6_submission.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_U4PLGH a_n321_n518# a_n33_118# a_15_549# a_207_n615#
+ a_n225_118# a_n413_118# a_111_21# a_n369_n615# a_207_549# a_n33_n518# a_111_n87#
+ a_63_118# a_15_n615# w_n551_n737# a_n177_n615# a_255_118# a_n177_549# a_159_n518#
+ a_n81_21# a_n273_21# a_303_21# a_n413_n518# a_303_n87# a_n129_118# a_255_n518# a_n369_549#
+ a_351_n518# a_n81_n87# a_n321_118# a_n273_n87# a_n129_n518# a_63_n518# a_159_118#
+ a_n225_n518# a_351_118#
X0 a_63_n518# a_15_n615# a_n33_n518# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n129_n518# a_n177_n615# a_n225_n518# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_n33_n518# a_n81_n87# a_n129_n518# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 a_351_n518# a_303_n87# a_255_n518# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n33_118# a_n81_21# a_n129_118# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_351_118# a_303_21# a_255_118# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_159_118# a_111_21# a_63_118# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_255_118# a_207_549# a_159_118# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 a_n321_118# a_n369_549# a_n413_118# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X9 a_n225_118# a_n273_21# a_n321_118# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X10 a_n129_118# a_n177_549# a_n225_118# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 a_255_n518# a_207_n615# a_159_n518# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_n321_n518# a_n369_n615# a_n413_n518# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X13 a_63_118# a_15_549# a_n33_118# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 a_159_n518# a_111_n87# a_63_n518# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 a_n225_n518# a_n273_n87# a_n321_n518# w_n551_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_PDCJZ5 a_n345_n200# a_29_n297# a_n129_n297# a_187_n297#
+ a_129_n200# a_n287_n297# a_287_n200# w_n483_n419# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n483_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_287_n200# a_187_n297# a_129_n200# w_n483_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2 a_129_n200# a_29_n297# a_n29_n200# w_n483_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3 a_n29_n200# a_n129_n297# a_n187_n200# w_n483_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
.ends

.subckt bias_curm_p m1_216_n466# m1_120_n692# a_172_n788# w_172_376#
Xsky130_fd_pr__pfet_01v8_U4PLGH_0 m1_216_n466# m1_120_n692# a_172_n788# a_172_n788#
+ m1_120_n692# m1_120_n692# a_172_n788# a_172_n788# a_172_n788# m1_120_n692# a_172_n788#
+ m1_216_n466# a_172_n788# w_172_376# a_172_n788# m1_216_n466# a_172_n788# m1_120_n692#
+ a_172_n788# a_172_n788# a_172_n788# m1_120_n692# a_172_n788# m1_216_n466# m1_216_n466#
+ a_172_n788# m1_120_n692# a_172_n788# m1_216_n466# a_172_n788# m1_216_n466# m1_216_n466#
+ m1_120_n692# m1_120_n692# m1_120_n692# sky130_fd_pr__pfet_01v8_U4PLGH
Xsky130_fd_pr__pfet_01v8_PDCJZ5_0 m1_120_n692# a_172_n788# a_172_n788# a_172_n788#
+ w_172_376# a_172_n788# m1_120_n692# w_172_376# m1_120_n692# w_172_376# sky130_fd_pr__pfet_01v8_PDCJZ5
.ends

.subckt curr_mirror_distribution m2_290_1950# I_in m3_1720_60#
Xbias_curm_p_6 I_out4 bias_curm_p_6/m1_120_n692# I_in m2_290_1950# bias_curm_p
Xbias_curm_p_7 I_out8 bias_curm_p_7/m1_120_n692# I_in m2_290_1950# bias_curm_p
Xbias_curm_p_8 I_out7 bias_curm_p_8/m1_120_n692# I_in m2_290_1950# bias_curm_p
Xbias_curm_p_0 I_in bias_curm_p_0/m1_120_n692# I_in m2_290_1950# bias_curm_p
Xbias_curm_p_1 m3_1720_60# bias_curm_p_1/m1_120_n692# I_in m2_290_1950# bias_curm_p
Xbias_curm_p_2 I_out2 bias_curm_p_2/m1_120_n692# I_in m2_290_1950# bias_curm_p
Xbias_curm_p_3 I_out3 bias_curm_p_3/m1_120_n692# I_in m2_290_1950# bias_curm_p
Xbias_curm_p_4 I_out6 bias_curm_p_4/m1_120_n692# I_in m2_290_1950# bias_curm_p
Xbias_curm_p_5 I_out5 bias_curm_p_5/m1_120_n692# I_in m2_290_1950# bias_curm_p
.ends

.subckt sky130_fd_pr__nfet_01v8_CDW43Z a_100_n50# a_n100_n138# a_n260_n224# a_n158_n50#
X0 a_100_n50# a_n100_n138# a_n158_n50# a_n260_n224# sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_F8VELN a_n513_n200# a_n129_n200# a_399_n288# a_63_n200#
+ a_n225_n200# a_495_222# a_111_222# a_n321_n200# a_207_n288# a_n33_n200# a_n369_n288#
+ a_n707_n374# a_303_222# a_n605_n200# a_447_n200# a_15_n288# a_n81_222# a_n177_n288#
+ a_n561_n288# a_543_n200# a_159_n200# a_n273_222# a_255_n200# a_351_n200# a_n417_n200#
+ a_n465_222#
X0 a_n33_n200# a_n81_222# a_n129_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_351_n200# a_303_222# a_255_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_255_n200# a_207_n288# a_159_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n321_n200# a_n369_n288# a_n417_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_543_n200# a_495_222# a_447_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_159_n200# a_111_222# a_63_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_n225_n200# a_n273_222# a_n321_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X7 a_447_n200# a_399_n288# a_351_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 a_n513_n200# a_n561_n288# a_n605_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X9 a_63_n200# a_15_n288# a_n33_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 a_n129_n200# a_n177_n288# a_n225_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 a_n417_n200# a_n465_222# a_n513_n200# a_n707_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_854667 a_n287_n200# a_745_n200# a_n487_n288# a_545_n288#
+ a_229_n200# a_n545_n200# a_29_n288# a_n745_n288# a_487_n200# a_n29_n200# a_n229_n288#
+ a_n905_n374# a_287_n288# a_n803_n200#
X0 a_745_n200# a_545_n288# a_487_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X1 a_487_n200# a_287_n288# a_229_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X2 a_n29_n200# a_n229_n288# a_n287_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X3 a_229_n200# a_29_n288# a_n29_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4 a_n545_n200# a_n745_n288# a_n803_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X5 a_n287_n200# a_n487_n288# a_n545_n200# a_n905_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
.ends

.subckt tia_cur_mirror m1_71_n690# a_122_42# m1_71_130# m1_167_370# VSUBS
Xsky130_fd_pr__nfet_01v8_F8VELN_0 m1_167_370# m1_167_370# a_122_42# m1_167_370# m1_71_130#
+ a_122_42# a_122_42# m1_167_370# a_122_42# m1_71_130# a_122_42# VSUBS a_122_42# m1_71_130#
+ m1_167_370# a_122_42# a_122_42# a_122_42# a_122_42# m1_71_130# m1_71_130# a_122_42#
+ m1_167_370# m1_71_130# m1_71_130# a_122_42# sky130_fd_pr__nfet_01v8_F8VELN
Xsky130_fd_pr__nfet_01v8_854667_0 m1_71_n690# m1_71_n690# a_122_42# a_122_42# m1_71_n690#
+ m1_71_130# a_122_42# a_122_42# m1_71_130# m1_71_130# a_122_42# VSUBS a_122_42# m1_71_n690#
+ sky130_fd_pr__nfet_01v8_854667
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ZRA4RB a_n523_21# a_n817_n597# a_n1156_n509# a_n523_n87#
+ a_n1209_531# a_608_n509# a_216_109# a_n862_n509# a_n621_n597# a_n1209_n597# a_n568_109#
+ a_n78_n509# a_706_109# a_653_21# a_412_n509# a_653_n87# a_n817_531# a_n327_21# a_n131_n87#
+ a_n78_109# a_n1254_n509# a_n1058_109# a_n1013_n597# a_706_n509# a_n176_109# a_359_n597#
+ a_314_109# a_n176_n509# a_947_531# a_261_n87# a_n960_n509# a_n425_531# a_1143_n597#
+ a_457_21# a_n1111_n87# a_510_n509# a_n666_109# a_804_109# a_65_21# a_163_n597# a_n229_n597#
+ a_n1356_n683# a_n1156_109# a_555_531# a_804_n509# a_n274_n509# a_n915_21# a_n274_109#
+ a_412_109# a_1098_n509# a_n719_n87# a_n33_n597# a_1098_109# a_163_531# a_n764_109#
+ a_902_109# a_n568_n509# a_n33_531# a_n131_21# a_n1013_531# a_118_n509# a_902_n509#
+ a_n1254_109# a_849_n87# a_n719_21# a_n327_n87# a_555_n597# a_n372_n509# a_n1111_21#
+ a_1196_n509# a_1143_531# a_n372_109# a_510_109# a_261_21# a_20_109# a_n621_531#
+ a_1196_109# a_n666_n509# a_1000_109# a_n425_n597# a_849_21# a_n862_109# a_457_n87#
+ a_216_n509# a_1000_n509# a_751_531# a_n470_n509# a_n1058_n509# a_118_109# a_n470_109#
+ a_n229_531# a_n915_n87# a_947_n597# a_n764_n509# a_20_n509# a_608_109# a_1045_21#
+ a_n960_109# a_314_n509# a_65_n87# a_359_531# a_751_n597# a_1045_n87#
X0 a_n274_109# a_n327_21# a_n372_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X1 a_n764_n509# a_n817_n597# a_n862_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X2 a_706_n509# a_653_n87# a_608_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X3 a_n568_109# a_n621_531# a_n666_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X4 a_n862_109# a_n915_21# a_n960_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X5 a_1196_n509# a_1143_n597# a_1098_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X6 a_1196_109# a_1143_531# a_1098_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X7 a_n1156_n509# a_n1209_n597# a_n1254_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X8 a_n960_109# a_n1013_531# a_n1058_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X9 a_412_109# a_359_531# a_314_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X10 a_n470_n509# a_n523_n87# a_n568_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X11 a_n372_n509# a_n425_n597# a_n470_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X12 a_314_n509# a_261_n87# a_216_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X13 a_706_109# a_653_21# a_608_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X14 a_n862_n509# a_n915_n87# a_n960_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X15 a_n78_109# a_n131_21# a_n176_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X16 a_1000_109# a_947_531# a_902_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X17 a_804_n509# a_751_n597# a_706_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X18 a_n372_109# a_n425_531# a_n470_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X19 a_118_n509# a_65_n87# a_20_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X20 a_n666_109# a_n719_21# a_n764_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X21 a_n78_n509# a_n131_n87# a_n176_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X22 a_n1058_109# a_n1111_21# a_n1156_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X23 a_n568_n509# a_n621_n597# a_n666_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X24 a_412_n509# a_359_n597# a_314_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X25 a_216_109# a_163_531# a_118_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X26 a_118_109# a_65_21# a_20_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X27 a_510_109# a_457_21# a_412_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X28 a_n960_n509# a_n1013_n597# a_n1058_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X29 a_902_n509# a_849_n87# a_804_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X30 a_804_109# a_751_531# a_706_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X31 a_n176_109# a_n229_531# a_n274_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X32 a_n176_n509# a_n229_n597# a_n274_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X33 a_n470_109# a_n523_21# a_n568_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X34 a_n764_109# a_n817_531# a_n862_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X35 a_n666_n509# a_n719_n87# a_n764_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X36 a_510_n509# a_457_n87# a_412_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X37 a_1098_109# a_1045_21# a_1000_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X38 a_608_n509# a_555_n597# a_510_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X39 a_20_109# a_n33_531# a_n78_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X40 a_n1156_109# a_n1209_531# a_n1254_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X41 a_1000_n509# a_947_n597# a_902_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X42 a_1098_n509# a_1045_n87# a_1000_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X43 a_314_109# a_261_21# a_216_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X44 a_n1058_n509# a_n1111_n87# a_n1156_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X45 a_608_109# a_555_531# a_510_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X46 a_n274_n509# a_n327_n87# a_n372_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X47 a_902_109# a_849_21# a_804_109# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X48 a_20_n509# a_n33_n597# a_n78_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X49 a_216_n509# a_163_n597# a_118_n509# a_n1356_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
.ends

.subckt sky130_fd_pr__pfet_01v8_NZHYX4 a_n568_n518# a_n764_118# a_653_n615# a_n719_n615#
+ a_163_n87# a_n33_n87# a_118_n518# a_n372_n518# a_n523_n615# a_510_118# a_n372_118#
+ a_20_118# a_65_549# a_n666_n518# a_n621_n87# a_163_21# a_n523_549# a_216_n518# a_n470_n518#
+ w_n902_n737# a_118_118# a_n470_118# a_653_549# a_n131_549# a_20_n518# a_n764_n518#
+ a_n229_n87# a_n621_21# a_314_n518# a_608_118# a_65_n615# a_359_n87# a_n33_21# a_261_549#
+ a_608_n518# a_216_118# a_n425_21# a_412_n518# a_n78_n518# a_706_118# a_n568_118#
+ a_457_n615# a_n78_118# a_555_21# a_n719_549# a_706_n518# a_n229_21# a_314_118# a_n176_118#
+ a_n176_n518# a_261_n615# a_n327_n615# a_510_n518# a_n425_n87# a_n666_118# a_359_21#
+ a_n327_549# a_n131_n615# a_n274_n518# a_555_n87# a_457_549# a_412_118# a_n274_118#
X0 a_n666_n518# a_n719_n615# a_n764_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X1 a_510_n518# a_457_n615# a_412_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X2 a_20_118# a_n33_21# a_n78_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X3 a_608_n518# a_555_n87# a_510_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X4 a_314_118# a_261_549# a_216_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X5 a_608_118# a_555_21# a_510_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X6 a_n274_n518# a_n327_n615# a_n372_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X7 a_20_n518# a_n33_n87# a_n78_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X8 a_216_n518# a_163_n87# a_118_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X9 a_n274_118# a_n327_549# a_n372_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X10 a_706_n518# a_653_n615# a_608_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X11 a_n568_118# a_n621_21# a_n666_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X12 a_412_118# a_359_21# a_314_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X13 a_n470_n518# a_n523_n615# a_n568_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X14 a_n372_n518# a_n425_n87# a_n470_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X15 a_314_n518# a_261_n615# a_216_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X16 a_706_118# a_653_549# a_608_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X17 a_n78_118# a_n131_549# a_n176_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X18 a_n372_118# a_n425_21# a_n470_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X19 a_118_n518# a_65_n615# a_20_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X20 a_n666_118# a_n719_549# a_n764_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X21 a_n78_n518# a_n131_n615# a_n176_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X22 a_n568_n518# a_n621_n87# a_n666_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X23 a_412_n518# a_359_n87# a_314_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X24 a_118_118# a_65_549# a_20_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X25 a_216_118# a_163_21# a_118_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X26 a_510_118# a_457_549# a_412_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X27 a_n176_118# a_n229_21# a_n274_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X28 a_n176_n518# a_n229_n87# a_n274_n518# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X29 a_n470_118# a_n523_549# a_n568_118# w_n902_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
.ends

.subckt rf_transistors m1_2957_359# m1_1943_755# m1_2041_n2774# m1_3839_995# m1_1257_995#
+ m1_1551_n2534# m1_2727_n2534# m1_3643_119# m1_1061_119# m1_1061_n1330# m1_865_995#
+ m1_2237_n1330# m1_571_n2534# m1_1453_n472# m1_1747_359# m1_2761_755# m1_1061_n1916#
+ m1_2237_n1916# m1_3021_n472# m1_767_n712# m1_669_119# m1_1943_n2156# m1_2139_n2534#
+ a_622_n800# m1_1649_n2774# m1_2565_359# m1_1551_755# m1_963_n2156# m1_3447_995#
+ m1_1943_n1090# m1_3251_119# m1_669_n2774# m1_963_n1090# m1_2825_n2774# m1_571_n712#
+ m1_669_n472# m1_1355_359# m1_1159_n712# m1_1845_n1330# m1_1355_n2156# m1_963_359#
+ m1_2041_119# m1_1943_n712# m1_2335_n712# m1_865_n1330# m1_1845_n1916# m1_2369_755#
+ m1_1355_n1090# m1_2531_n2156# m1_3741_755# m1_3055_995# m1_865_n1916# m1_1061_n2774#
+ m1_2237_n2774# m1_2531_n1090# m1_1747_n2534# m1_2859_119# m1_1845_995# m1_1257_n1330#
+ m1_3545_359# m1_1159_755# m1_767_n2534# m1_1845_n472# m1_2237_n472# m1_2923_n2534#
+ m1_767_755# m1_571_359# m1_1257_n1916# a_623_n2862# m1_2433_n1330# m1_1649_119#
+ m1_2663_995# a_622_n2244# m1_2433_n1916# m1_1159_n2534# m1_2467_119# m1_1453_995#
+ m1_2335_n2534# m1_2041_n472# m1_3349_755# a_623_658# m1_1845_n2774# m1_3153_359#
+ m1_963_n712# m1_1943_359# m1_865_n2774# m1_3839_119# m1_1257_119# m1_3021_n1330#
+ m1_865_119# m1_2727_n712# m1_1551_n2156# m1_2727_n2156# m1_2957_755# m1_2761_359#
+ m1_3021_n1916# m1_3643_995# m1_571_n2156# m1_1257_n2774# a_623_22# m1_1061_995#
+ m1_1551_n1090# m1_2727_n1090# m1_865_n472# m1_1355_n712# m1_2433_n2774# m1_1747_755#
+ m1_571_n1090# m1_1943_n2534# m1_1551_359# m1_2629_n472# m1_2531_n712# m1_3447_119#
+ m1_1453_n1330# m1_2629_n1330# m1_2139_n2156# m1_669_995# m1_963_n2534# w_623_22#
+ m1_1453_n1916# m1_2565_755# m1_2139_n1090# m1_2629_n1916# m1_1257_n472# m1_3251_995#
+ a_623_n908# a_2421_658# m1_2433_n472# m1_1355_n2534# m1_2369_359# m1_3741_359# m1_1355_755#
+ m1_3021_n2774# m1_3055_119# m1_963_755# m1_2041_995# m1_2531_n2534# a_2421_22# m1_2041_n1330#
+ m1_1845_119# m1_1061_n472# m1_1159_359# m1_1747_n2156# m1_767_359# m1_2041_n1916#
+ m1_2859_995# m1_767_n2156# m1_1747_n1090# m1_2923_n2156# m1_2663_119# m1_3545_755#
+ m1_1747_n712# m1_1453_n2774# m1_2139_n712# m1_767_n1090# m1_2629_n2774# m1_571_755#
+ m1_2923_n712# m1_2923_n1090# m1_1649_995# m1_1649_n1330# m1_1159_n2156# m1_1453_119#
+ m1_3349_359# m1_669_n1330# m1_1649_n1916# m1_1159_n1090# m1_2825_n1330# m1_2335_n2156#
+ m1_1551_n712# m1_1649_n472# m1_2467_995# m1_669_n1916# m1_3153_755# VSUBS m1_2825_n472#
+ m1_2335_n1090# m1_2825_n1916#
Xsky130_fd_pr__nfet_01v8_lvt_ZRA4RB_0 a_622_n2244# a_623_n2862# m1_669_n2774# a_623_n2862#
+ a_622_n2244# m1_2433_n2774# m1_2041_n1916# m1_963_n2534# a_623_n2862# a_623_n2862#
+ m1_1257_n1916# m1_1747_n2534# m1_2531_n2156# a_622_n2244# m1_2237_n2774# a_623_n2862#
+ a_622_n2244# a_622_n2244# a_623_n2862# m1_1747_n2156# m1_571_n2534# m1_767_n2156#
+ a_623_n2862# m1_2531_n2534# m1_1649_n1916# a_623_n2862# m1_2139_n2156# m1_1649_n2774#
+ a_622_n2244# a_623_n2862# m1_865_n2774# a_622_n2244# a_623_n2862# a_622_n2244# a_623_n2862#
+ m1_2335_n2534# m1_1159_n2156# m1_2629_n1916# a_622_n2244# a_623_n2862# a_623_n2862#
+ VSUBS m1_669_n1916# a_622_n2244# m1_2629_n2774# m1_1551_n2534# a_622_n2244# m1_1551_n2156#
+ m1_2237_n1916# m1_2923_n2534# a_623_n2862# a_623_n2862# m1_2923_n2156# a_622_n2244#
+ m1_1061_n1916# m1_2727_n2156# m1_1257_n2774# a_622_n2244# a_622_n2244# a_622_n2244#
+ m1_1943_n2534# m1_2727_n2534# m1_571_n2156# a_623_n2862# a_622_n2244# a_623_n2862#
+ a_623_n2862# m1_1453_n2774# a_622_n2244# m1_3021_n2774# a_622_n2244# m1_1453_n1916#
+ m1_2335_n2156# a_622_n2244# m1_1845_n1916# a_622_n2244# m1_3021_n1916# m1_1159_n2534#
+ m1_2825_n1916# a_623_n2862# a_622_n2244# m1_963_n2156# a_623_n2862# m1_2041_n2774#
+ m1_2825_n2774# a_622_n2244# m1_1355_n2534# m1_767_n2534# m1_1943_n2156# m1_1355_n2156#
+ a_622_n2244# a_623_n2862# a_623_n2862# m1_1061_n2774# m1_1845_n2774# m1_2433_n1916#
+ a_622_n2244# m1_865_n1916# m1_2139_n2534# a_623_n2862# a_622_n2244# a_623_n2862#
+ a_623_n2862# sky130_fd_pr__nfet_01v8_lvt_ZRA4RB
Xsky130_fd_pr__nfet_01v8_lvt_ZRA4RB_1 a_622_n800# a_623_n908# m1_669_n1330# a_623_n908#
+ a_622_n800# m1_2433_n1330# m1_2041_n472# m1_963_n1090# a_623_n908# a_623_n908# m1_1257_n472#
+ m1_1747_n1090# m1_2531_n712# a_622_n800# m1_2237_n1330# a_623_n908# a_622_n800#
+ a_622_n800# a_623_n908# m1_1747_n712# m1_571_n1090# m1_767_n712# a_623_n908# m1_2531_n1090#
+ m1_1649_n472# a_623_n908# m1_2139_n712# m1_1649_n1330# a_622_n800# a_623_n908# m1_865_n1330#
+ a_622_n800# a_623_n908# a_622_n800# a_623_n908# m1_2335_n1090# m1_1159_n712# m1_2629_n472#
+ a_622_n800# a_623_n908# a_623_n908# VSUBS m1_669_n472# a_622_n800# m1_2629_n1330#
+ m1_1551_n1090# a_622_n800# m1_1551_n712# m1_2237_n472# m1_2923_n1090# a_623_n908#
+ a_623_n908# m1_2923_n712# a_622_n800# m1_1061_n472# m1_2727_n712# m1_1257_n1330#
+ a_622_n800# a_622_n800# a_622_n800# m1_1943_n1090# m1_2727_n1090# m1_571_n712# a_623_n908#
+ a_622_n800# a_623_n908# a_623_n908# m1_1453_n1330# a_622_n800# m1_3021_n1330# a_622_n800#
+ m1_1453_n472# m1_2335_n712# a_622_n800# m1_1845_n472# a_622_n800# m1_3021_n472#
+ m1_1159_n1090# m1_2825_n472# a_623_n908# a_622_n800# m1_963_n712# a_623_n908# m1_2041_n1330#
+ m1_2825_n1330# a_622_n800# m1_1355_n1090# m1_767_n1090# m1_1943_n712# m1_1355_n712#
+ a_622_n800# a_623_n908# a_623_n908# m1_1061_n1330# m1_1845_n1330# m1_2433_n472#
+ a_622_n800# m1_865_n472# m1_2139_n1090# a_623_n908# a_622_n800# a_623_n908# a_623_n908#
+ sky130_fd_pr__nfet_01v8_lvt_ZRA4RB
Xsky130_fd_pr__pfet_01v8_NZHYX4_1 m1_767_359# m1_571_755# a_623_22# a_623_22# a_623_22#
+ a_623_22# m1_1453_119# m1_963_359# a_623_22# m1_1845_995# m1_963_755# m1_1355_755#
+ a_623_658# m1_669_119# a_623_22# a_623_658# a_623_658# m1_1551_359# m1_865_119#
+ w_623_22# m1_1453_995# m1_865_995# a_623_658# a_623_658# m1_1355_359# m1_571_359#
+ a_623_22# a_623_658# m1_1649_119# m1_1943_755# a_623_22# a_623_22# a_623_658# a_623_658#
+ m1_1943_359# m1_1551_755# a_623_658# m1_1747_359# m1_1257_119# m1_2041_995# m1_767_755#
+ a_623_22# m1_1257_995# a_623_658# a_623_658# m1_2041_119# a_623_658# m1_1649_995#
+ m1_1159_755# m1_1159_359# a_623_22# a_623_22# m1_1845_119# a_623_22# m1_669_995#
+ a_623_658# a_623_658# a_623_22# m1_1061_119# a_623_22# a_623_658# m1_1747_755# m1_1061_995#
+ sky130_fd_pr__pfet_01v8_NZHYX4
Xsky130_fd_pr__pfet_01v8_NZHYX4_2 m1_2565_359# m1_2369_755# a_2421_22# a_2421_22#
+ a_2421_22# a_2421_22# m1_3251_119# m1_2761_359# a_2421_22# m1_3643_995# m1_2761_755#
+ m1_3153_755# a_2421_658# m1_2467_119# a_2421_22# a_2421_658# a_2421_658# m1_3349_359#
+ m1_2663_119# w_623_22# m1_3251_995# m1_2663_995# a_2421_658# a_2421_658# m1_3153_359#
+ m1_2369_359# a_2421_22# a_2421_658# m1_3447_119# m1_3741_755# a_2421_22# a_2421_22#
+ a_2421_658# a_2421_658# m1_3741_359# m1_3349_755# a_2421_658# m1_3545_359# m1_3055_119#
+ m1_3839_995# m1_2565_755# a_2421_22# m1_3055_995# a_2421_658# a_2421_658# m1_3839_119#
+ a_2421_658# m1_3447_995# m1_2957_755# m1_2957_359# a_2421_22# a_2421_22# m1_3643_119#
+ a_2421_22# m1_2467_995# a_2421_658# a_2421_658# a_2421_22# m1_2859_119# a_2421_22#
+ a_2421_658# m1_3545_755# m1_2859_995# sky130_fd_pr__pfet_01v8_NZHYX4
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_ZWVPUJ m4_n2851_n1900# c2_n2751_n1800#
X0 c2_n2751_n1800# m4_n2851_n1900# sky130_fd_pr__cap_mim_m3_2 l=1.8e+07u w=2.5e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_RRWALQ a_n1041_109# a_n1041_727# a_1119_1149# a_n1185_21#
+ a_n1229_109# a_n1229_727# a_n753_n509# a_879_n1127# a_n81_727# a_447_639# a_n369_n509#
+ a_687_n1127# a_975_n1127# a_n81_109# a_n129_531# a_351_n87# a_399_n1127# a_495_n1127#
+ a_783_n1127# a_n33_n87# a_399_727# a_303_n509# a_591_n1127# a_399_109# a_n513_n597#
+ a_n129_n597# a_n321_639# a_879_109# a_879_727# a_63_n597# a_n273_109# a_n273_727#
+ a_n1089_n597# a_735_21# a_447_531# a_n225_n87# a_n465_n509# a_n753_727# a_n753_109#
+ a_n225_1149# a_15_109# a_15_727# a_n705_n705# a_1167_n509# a_255_n705# a_n321_531#
+ a_927_1149# a_n1185_1149# a_591_109# a_591_727# a_15_n509# a_n609_21# a_1119_21#
+ a_639_639# a_543_n87# a_n561_n509# a_1071_109# a_1071_727# a_1119_n1215# a_n177_n509#
+ a_n993_21# a_n33_n1215# a_207_727# a_n897_639# a_n321_n597# a_111_n509# a_207_109#
+ a_879_n509# a_n513_639# a_n609_n1215# a_n417_n1215# a_n1229_n1127# a_n465_727# a_639_n597#
+ a_n1185_n1215# a_n465_109# a_1023_n597# a_n801_n1215# a_n225_n1215# a_639_531# a_n417_n87#
+ a_n1137_n509# a_n273_n509# a_351_21# a_n945_727# a_n945_109# a_n1331_n1301# a_n897_531#
+ a_975_n509# a_831_639# a_n513_531# a_n513_n705# a_n129_n705# a_735_1149# a_n33_1149#
+ a_783_727# a_927_n1215# a_783_109# a_735_n1215# a_159_n1215# a_735_n87# a_543_n1215#
+ a_n33_21# a_n225_21# a_63_n705# a_351_n1215# a_n1089_n705# a_927_21# a_n1089_639#
+ a_15_n1127# a_n993_n87# a_n177_727# a_n177_109# a_831_531# a_n705_639# a_687_n509#
+ a_n897_n597# a_1071_n509# a_n657_727# a_831_n597# a_n657_109# a_447_n597# a_n993_n1215#
+ a_n609_n87# a_n1137_727# a_n1137_109# a_1023_639# a_n1089_531# a_495_727# a_n993_1149#
+ a_495_109# a_n1137_n1127# a_n705_531# a_111_727# a_n81_n509# a_783_n509# a_111_109#
+ a_n849_n509# a_399_n509# a_n321_n705# a_n1041_n1127# a_975_727# a_543_1149# a_63_639#
+ a_975_109# a_n609_1149# a_159_1149# a_927_n87# a_639_n705# a_n1041_n509# a_1023_n705#
+ a_1023_531# a_n1185_n87# a_543_21# a_n369_727# a_n369_109# a_159_21# a_n801_n87#
+ a_n945_n509# a_495_n509# a_207_n1127# a_n849_109# a_63_531# a_n849_727# a_255_639#
+ a_303_n1127# a_111_n1127# a_n705_n597# a_255_n597# a_1167_n1127# a_n801_21# a_159_n87#
+ a_n81_n1127# a_n417_21# a_1071_n1127# a_687_727# a_n1229_n509# a_687_109# a_303_727#
+ a_n849_n1127# a_303_109# a_1167_727# a_591_n509# a_1167_109# a_n657_n509# a_n945_n1127#
+ a_n657_n1127# a_n369_n1127# a_n897_n705# a_255_531# a_n129_639# a_n801_1149# a_1119_n87#
+ a_n753_n1127# a_n465_n1127# a_n177_n1127# a_351_1149# a_n561_n1127# a_n561_727#
+ a_n417_1149# a_n273_n1127# a_n561_109# a_831_n705# a_207_n509# a_447_n705#
X0 a_111_727# a_63_639# a_15_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_15_109# a_n33_21# a_n81_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_1071_n509# a_1023_n597# a_975_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n81_727# a_n129_639# a_n177_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n273_727# a_n321_639# a_n369_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_n177_727# a_n225_1149# a_n273_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 a_399_n509# a_351_n87# a_303_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_399_n1127# a_351_n1215# a_303_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X8 a_111_109# a_63_531# a_15_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X9 a_n465_n509# a_n513_n597# a_n561_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_n81_109# a_n129_531# a_n177_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X11 a_879_n1127# a_831_n705# a_783_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_n273_109# a_n321_531# a_n369_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X13 a_687_n509# a_639_n597# a_591_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X14 a_1071_n1127# a_1023_n705# a_975_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X15 a_n177_109# a_n225_21# a_n273_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 a_n81_n1127# a_n129_n705# a_n177_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17 a_n753_n509# a_n801_n87# a_n849_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X18 a_495_n1127# a_447_n705# a_399_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X19 a_n657_n1127# a_n705_n705# a_n753_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X20 a_975_n509# a_927_n87# a_879_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X21 a_975_n1127# a_927_n1215# a_879_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 a_n1137_n1127# a_n1185_n1215# a_n1229_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X23 a_n81_n509# a_n129_n597# a_n177_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X24 a_15_n509# a_n33_n87# a_n81_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X25 a_591_n1127# a_543_n1215# a_495_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X26 a_n753_n1127# a_n801_n1215# a_n849_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X27 a_n369_n509# a_n417_n87# a_n465_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X28 a_n1041_n509# a_n1089_n597# a_n1137_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X29 a_15_n1127# a_n33_n1215# a_n81_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X30 a_n657_n509# a_n705_n597# a_n753_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X31 a_879_n509# a_831_n597# a_783_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X32 a_n945_n509# a_n993_n87# a_n1041_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X33 a_1167_n509# a_1119_n87# a_1071_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X34 a_1167_n1127# a_1119_n1215# a_1071_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X35 a_n177_n1127# a_n225_n1215# a_n273_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X36 a_303_n509# a_255_n597# a_207_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X37 a_n273_n509# a_n321_n597# a_n369_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X38 a_303_727# a_255_639# a_207_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X39 a_591_727# a_543_1149# a_495_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X40 a_591_n509# a_543_n87# a_495_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X41 a_783_727# a_735_1149# a_687_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X42 a_495_727# a_447_639# a_399_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X43 a_207_727# a_159_1149# a_111_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 a_207_n1127# a_159_n1215# a_111_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X45 a_111_n1127# a_63_n705# a_15_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 a_n273_n1127# a_n321_n705# a_n369_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X47 a_975_727# a_927_1149# a_879_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X48 a_687_727# a_639_639# a_591_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 a_399_727# a_351_1149# a_303_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 a_n369_n1127# a_n417_n1215# a_n465_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X51 a_879_727# a_831_639# a_783_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 a_687_n1127# a_639_n705# a_591_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X53 a_n1041_727# a_n1089_639# a_n1137_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X54 a_n849_n1127# a_n897_n705# a_n945_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X55 a_n1137_727# a_n1185_1149# a_n1229_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X56 a_n849_n509# a_n897_n597# a_n945_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X57 a_1071_727# a_1023_639# a_975_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X58 a_n561_727# a_n609_1149# a_n657_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X59 a_303_n1127# a_255_n705# a_207_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 a_1167_727# a_1119_1149# a_1071_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X61 a_n465_727# a_n513_639# a_n561_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X62 a_n753_727# a_n801_1149# a_n849_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X63 a_n945_727# a_n993_1149# a_n1041_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X64 a_207_n509# a_159_n87# a_111_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X65 a_591_109# a_543_21# a_495_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X66 a_303_109# a_255_531# a_207_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X67 a_n369_727# a_n417_1149# a_n465_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 a_n657_727# a_n705_639# a_n753_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X69 a_n465_n1127# a_n513_n705# a_n561_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X70 a_207_109# a_159_21# a_111_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 a_n849_727# a_n897_639# a_n945_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X72 a_783_n1127# a_735_n1215# a_687_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 a_n177_n509# a_n225_n87# a_n273_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 a_783_109# a_735_21# a_687_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X75 a_495_109# a_447_531# a_399_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X76 a_687_109# a_639_531# a_591_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X77 a_399_109# a_351_21# a_303_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 a_975_109# a_927_21# a_879_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X79 a_n945_n1127# a_n993_n1215# a_n1041_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X80 a_879_109# a_831_531# a_783_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 a_n1041_109# a_n1089_531# a_n1137_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X82 a_15_727# a_n33_1149# a_n81_727# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X83 a_495_n509# a_447_n597# a_399_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 a_n1137_109# a_n1185_21# a_n1229_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X85 a_n1137_n509# a_n1185_n87# a_n1229_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X86 a_1071_109# a_1023_531# a_975_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X87 a_n561_n1127# a_n609_n1215# a_n657_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 a_n1041_n1127# a_n1089_n705# a_n1137_n1127# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 a_n561_109# a_n609_21# a_n657_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X90 a_n561_n509# a_n609_n87# a_n657_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 a_1167_109# a_1119_21# a_1071_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X92 a_n465_109# a_n513_531# a_n561_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X93 a_n753_109# a_n801_21# a_n849_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X94 a_111_n509# a_63_n597# a_15_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 a_n369_109# a_n417_21# a_n465_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 a_n657_109# a_n705_531# a_n753_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 a_n945_109# a_n993_21# a_n1041_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X98 a_783_n509# a_735_n87# a_687_n509# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X99 a_n849_109# a_n897_531# a_n945_109# a_n1331_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt dis_tran m1_1422_1633# m1_1038_1633# m1_174_1015# m1_2190_775# m1_1326_157#
+ m1_78_2011# m1_750_1393# m1_1806_775# m1_558_157# m1_366_1393# m1_462_2011# m1_2094_1015#
+ m1_1422_397# m1_270_1633# m1_1134_1015# m1_654_397# m1_2286_1393# m1_1710_1393#
+ m1_2382_2011# m1_1326_1393# m1_270_775# m1_1422_2011# m1_1038_775# m1_1038_2011#
+ m1_2190_1633# m1_942_2251# m1_750_157# m1_558_2251# m1_1230_1633# m1_1518_157# m1_1998_1633#
+ m1_2382_775# m1_174_1393# m1_1998_397# m1_2478_2251# m1_270_2011# m1_78_775# m1_1614_397#
+ m1_1902_2251# m1_1518_2251# m1_846_397# m1_90_1210# m1_1230_775# m1_2094_1393# m1_846_1633#
+ m1_1134_1393# m1_462_775# m1_2190_2011# m1_1710_157# m1_90_1830# m1_1230_2011# m1_2094_157#
+ m1_1998_2011# m1_942_157# m1_750_2251# m1_366_2251# m1_1806_1633# m1_942_1015# m1_2190_397#
+ m1_558_1015# m1_1806_397# m1_90_590# m1_2286_2251# m1_1710_2251# m1_1326_2251# m1_1422_775#
+ m1_174_157# m1_846_2011# m1_2478_1015# m1_90_2440# m1_654_775# m1_1902_1015# m1_1902_157#
+ m1_654_1633# m1_1518_1015# m1_2286_157# m1_270_397# m1_1038_397# m1_174_2251# m1_1806_2011#
+ m1_2382_397# m1_1614_1633# m1_750_1015# m1_366_1015# m1_1134_157# m1_2094_2251#
+ m1_942_1393# m1_1998_775# m1_558_1393# m1_78_1633# m1_1614_775# m1_78_397# m1_1134_2251#
+ m1_366_157# m1_654_2011# m1_2286_1015# m1_846_775# m1_90_70# m1_1710_1015# m1_1230_397#
+ m1_462_1633# m1_2478_157# m1_1326_1015# m1_2478_1393# m1_462_397# m1_1902_1393#
+ m1_1518_1393# m1_1614_2011# m1_2382_1633# VSUBS
Xsky130_fd_pr__nfet_01v8_RRWALQ_0 m1_270_1633# m1_270_2011# m1_90_2440# m1_90_1210#
+ m1_78_1633# m1_78_2011# m1_558_1015# m1_2190_397# m1_1230_2011# m1_90_1830# m1_942_1015#
+ m1_1998_397# m1_2286_157# m1_1230_1633# m1_90_1830# m1_90_1210# m1_1710_157# m1_1806_397#
+ m1_2094_157# m1_90_1210# m1_1710_2251# m1_1614_775# m1_1902_157# m1_1710_1393# m1_90_590#
+ m1_90_590# m1_90_1830# m1_2190_1633# m1_2190_2011# m1_90_590# m1_1038_1633# m1_1038_2011#
+ m1_90_590# m1_90_1210# m1_90_1830# m1_90_1210# m1_846_775# m1_558_2251# m1_558_1393#
+ m1_90_2440# m1_1326_1393# m1_1326_2251# m1_90_590# m1_2478_1015# m1_90_590# m1_90_1830#
+ m1_90_2440# m1_90_2440# m1_1902_1393# m1_1902_2251# m1_1326_1015# m1_90_1210# m1_90_1210#
+ m1_90_1830# m1_90_1210# m1_750_1015# m1_2382_1633# m1_2382_2011# m1_90_70# m1_1134_1015#
+ m1_90_1210# m1_90_70# m1_1518_2251# m1_90_1830# m1_90_590# m1_1422_775# m1_1518_1393#
+ m1_2190_775# m1_90_1830# m1_90_70# m1_90_70# m1_78_397# m1_846_2011# m1_90_590#
+ m1_90_70# m1_846_1633# m1_90_590# m1_90_70# m1_90_70# m1_90_1830# m1_90_1210# m1_174_1015#
+ m1_1038_775# m1_90_1210# m1_366_2251# m1_366_1393# VSUBS m1_90_1830# m1_2286_1015#
+ m1_90_1830# m1_90_1830# m1_90_590# m1_90_590# m1_90_2440# m1_90_2440# m1_2094_2251#
+ m1_90_70# m1_2094_1393# m1_90_70# m1_90_70# m1_90_1210# m1_90_70# m1_90_1210# m1_90_1210#
+ m1_90_590# m1_90_70# m1_90_590# m1_90_1210# m1_90_1830# m1_1326_157# m1_90_1210#
+ m1_1134_2251# m1_1134_1393# m1_90_1830# m1_90_1830# m1_1998_775# m1_90_590# m1_2382_775#
+ m1_654_2011# m1_90_590# m1_654_1633# m1_90_590# m1_90_70# m1_90_1210# m1_174_2251#
+ m1_174_1393# m1_90_1830# m1_90_1830# m1_1806_2011# m1_90_2440# m1_1806_1633# m1_174_157#
+ m1_90_1830# m1_1422_2011# m1_1230_775# m1_2094_1015# m1_1422_1633# m1_462_775# m1_1710_1015#
+ m1_90_590# m1_270_397# m1_2286_2251# m1_90_2440# m1_90_1830# m1_2286_1393# m1_90_2440#
+ m1_90_2440# m1_90_1210# m1_90_590# m1_270_775# m1_90_590# m1_90_1830# m1_90_1210#
+ m1_90_1210# m1_942_2251# m1_942_1393# m1_90_1210# m1_90_1210# m1_366_1015# m1_1806_775#
+ m1_1518_157# m1_462_1633# m1_90_1830# m1_462_2011# m1_90_1830# m1_1614_397# m1_1422_397#
+ m1_90_590# m1_90_590# m1_2478_157# m1_90_1210# m1_90_1210# m1_1230_397# m1_90_1210#
+ m1_2382_397# m1_1998_2011# m1_78_775# m1_1998_1633# m1_1614_2011# m1_462_397# m1_1614_1633#
+ m1_2478_2251# m1_1902_1015# m1_2478_1393# m1_654_775# m1_366_157# m1_654_397# m1_942_157#
+ m1_90_590# m1_90_1830# m1_90_1830# m1_90_2440# m1_90_1210# m1_558_157# m1_846_397#
+ m1_1134_157# m1_90_2440# m1_750_157# m1_750_2251# m1_90_2440# m1_1038_397# m1_750_1393#
+ m1_90_590# m1_1518_1015# m1_90_590# sky130_fd_pr__nfet_01v8_RRWALQ
.ends

.subckt sky130_fd_pr__pfet_01v8_GYVK57 a_n819_n200# a_n345_n200# a_29_n297# a_n129_n297#
+ a_187_n297# a_129_n200# a_n503_n200# a_n287_n297# a_345_n297# a_287_n200# a_n661_n200#
+ a_n445_n297# a_503_n297# a_445_n200# a_n603_n297# a_661_n297# w_n957_n419# a_603_n200#
+ a_n761_n297# a_761_n200# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_761_n200# a_661_n297# a_603_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2 a_287_n200# a_187_n297# a_129_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3 a_n345_n200# a_n445_n297# a_n503_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X4 a_129_n200# a_29_n297# a_n29_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X5 a_445_n200# a_345_n297# a_287_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X6 a_n503_n200# a_n603_n297# a_n661_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X7 a_n29_n200# a_n129_n297# a_n187_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X8 a_603_n200# a_503_n297# a_445_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X9 a_n661_n200# a_n761_n297# a_n819_n200# w_n957_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_62U3RB a_608_n509# a_216_109# a_163_n87# a_n33_n87#
+ a_n327_531# a_n866_n683# a_n78_n509# a_n568_109# a_412_n509# a_706_109# a_n78_109#
+ a_457_531# a_706_n509# a_65_n597# a_n621_n87# a_n176_n509# a_314_109# a_n176_109#
+ a_163_21# a_510_n509# a_n666_109# a_n229_n87# a_n621_21# a_n274_n509# a_457_n597#
+ a_412_109# a_n274_109# a_65_531# a_n523_531# a_359_n87# a_n33_21# a_n568_n509# a_261_n597#
+ a_n327_n597# a_n764_109# a_118_n509# a_n425_21# a_653_531# a_n131_531# a_n372_n509#
+ a_n131_n597# a_510_109# a_n372_109# a_20_109# a_555_21# a_n666_n509# a_261_531#
+ a_n229_21# a_216_n509# a_653_n597# a_n470_n509# a_n425_n87# a_n719_n597# a_118_109#
+ a_n470_109# a_359_21# a_20_n509# a_n764_n509# a_n523_n597# a_608_109# a_314_n509#
+ a_555_n87# a_n719_531#
X0 a_n274_109# a_n327_531# a_n372_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X1 a_706_n509# a_653_n597# a_608_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X2 a_n568_109# a_n621_21# a_n666_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X3 a_412_109# a_359_21# a_314_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X4 a_n470_n509# a_n523_n597# a_n568_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X5 a_n372_n509# a_n425_n87# a_n470_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X6 a_314_n509# a_261_n597# a_216_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X7 a_706_109# a_653_531# a_608_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X8 a_n78_109# a_n131_531# a_n176_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X9 a_n372_109# a_n425_21# a_n470_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X10 a_118_n509# a_65_n597# a_20_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X11 a_n666_109# a_n719_531# a_n764_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X12 a_n78_n509# a_n131_n597# a_n176_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X13 a_n568_n509# a_n621_n87# a_n666_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X14 a_412_n509# a_359_n87# a_314_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X15 a_216_109# a_163_21# a_118_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X16 a_118_109# a_65_531# a_20_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X17 a_510_109# a_457_531# a_412_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X18 a_n176_109# a_n229_21# a_n274_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X19 a_n176_n509# a_n229_n87# a_n274_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X20 a_n470_109# a_n523_531# a_n568_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X21 a_n666_n509# a_n719_n597# a_n764_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=200000u
X22 a_510_n509# a_457_n597# a_412_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=200000u
X23 a_608_n509# a_555_n87# a_510_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X24 a_20_109# a_n33_21# a_n78_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X25 a_314_109# a_261_531# a_216_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X26 a_608_109# a_555_21# a_510_109# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X27 a_n274_n509# a_n327_n597# a_n372_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X28 a_20_n509# a_n33_n87# a_n78_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X29 a_216_n509# a_163_n87# a_118_n509# a_n866_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
.ends

.subckt fb_transistor m1_6753_3028# m1_6285_4403# sky130_fd_pr__pfet_01v8_GYVK57_0/a_503_n297#
+ m1_6459_2410# m1_7145_3028# m1_5871_3268# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n761_n297#
+ m1_6263_3268# m1_7145_2650# m1_6753_2650# m1_6917_4403# m1_6263_2410# m1_5871_2410#
+ m1_7233_4403# w_5706_2166# sky130_fd_pr__pfet_01v8_GYVK57_0/a_661_n297# m1_6127_4163#
+ a_5923_2832# m1_6759_4163# m1_5969_3028# m1_7075_4163# sky130_fd_pr__pfet_01v8_GYVK57_0/a_29_n297#
+ m1_5969_2650# m1_6655_3268# m1_6601_4403# m1_7047_3268# m1_6165_3028# m1_7047_2410#
+ m1_6655_2410# m1_7341_3028# m1_6165_2650# m1_6443_4163# m1_7341_2650# m1_7391_4163#
+ sky130_fd_pr__pfet_01v8_GYVK57_0/a_n129_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n287_n297#
+ m1_5811_4163# m1_6557_3028# m1_6851_3268# m1_6067_3268# sky130_fd_pr__pfet_01v8_GYVK57_0/a_187_n297#
+ m1_6557_2650# m1_7243_3268# m1_6067_2410# m1_6361_3028# a_5923_3450# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n445_n297#
+ m1_7243_2410# m1_6851_2410# m1_6361_2650# sky130_fd_pr__pfet_01v8_GYVK57_0/a_345_n297#
+ m1_6949_3028# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n603_n297# m1_6949_2650# m1_6459_3268#
+ m1_5969_4403# dw_5500_1960#
Xsky130_fd_pr__pfet_01v8_GYVK57_0 m1_5811_4163# m1_6285_4403# sky130_fd_pr__pfet_01v8_GYVK57_0/a_29_n297#
+ sky130_fd_pr__pfet_01v8_GYVK57_0/a_n129_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_187_n297#
+ m1_6759_4163# m1_6127_4163# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n287_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_345_n297#
+ m1_6917_4403# m1_5969_4403# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n445_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_503_n297#
+ m1_7075_4163# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n603_n297# sky130_fd_pr__pfet_01v8_GYVK57_0/a_661_n297#
+ dw_5500_1960# m1_7233_4403# sky130_fd_pr__pfet_01v8_GYVK57_0/a_n761_n297# m1_7391_4163#
+ m1_6601_4403# m1_6443_4163# sky130_fd_pr__pfet_01v8_GYVK57
Xsky130_fd_pr__nfet_01v8_lvt_62U3RB_0 m1_7243_2410# m1_6851_3268# a_5923_2832# a_5923_2832#
+ a_5923_3450# w_5706_2166# m1_6557_2650# m1_6067_3268# m1_7047_2410# m1_7341_3028#
+ m1_6557_3028# a_5923_3450# m1_7341_2650# a_5923_2832# a_5923_2832# m1_6459_2410#
+ m1_6949_3028# m1_6459_3268# a_5923_3450# m1_7145_2650# m1_5969_3028# a_5923_2832#
+ a_5923_3450# m1_6361_2650# a_5923_2832# m1_7047_3268# m1_6361_3028# a_5923_3450#
+ a_5923_3450# a_5923_2832# a_5923_3450# m1_6067_2410# a_5923_2832# a_5923_2832# m1_5871_3268#
+ m1_6753_2650# a_5923_3450# a_5923_3450# a_5923_3450# m1_6263_2410# a_5923_2832#
+ m1_7145_3028# m1_6263_3268# m1_6655_3268# a_5923_3450# m1_5969_2650# a_5923_3450#
+ a_5923_3450# m1_6851_2410# a_5923_2832# m1_6165_2650# a_5923_2832# a_5923_2832#
+ m1_6753_3028# m1_6165_3028# a_5923_3450# m1_6655_2410# m1_5871_2410# a_5923_2832#
+ m1_7243_3268# m1_6949_2650# a_5923_2832# a_5923_3450# sky130_fd_pr__nfet_01v8_lvt_62U3RB
.ends

.subckt tia_one_tia m1_n1960_n3240# m1_1850_2290# m2_1800_2380# tia_cur_mirror_0/m1_71_130#
+ w_1686_386# w_1650_2620# tia_cur_mirror_0/a_122_42# m2_n1840_n2910# VSUBS m1_1540_1550#
Xtia_cur_mirror_0 VSUBS tia_cur_mirror_0/a_122_42# tia_cur_mirror_0/m1_71_130# w_1686_386#
+ VSUBS tia_cur_mirror
Xrf_transistors_0 m1_1540_1550# m1_1540_1550# m2_n1840_n2910# w_1650_2620# w_1650_2620#
+ m1_1540_1550# m1_1540_1550# w_1650_2620# w_1650_2620# m2_n1840_n2910# w_1650_2620#
+ m2_n1840_n2910# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m2_n1840_n2910#
+ m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550# w_1650_2620# m1_1540_1550# m1_1540_1550#
+ w_1686_386# m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m1_1540_1550# w_1650_2620#
+ m1_1540_1550# w_1650_2620# m2_n1840_n2910# m1_1540_1550# m2_n1840_n2910# m1_1540_1550#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# m1_1540_1550#
+ w_1650_2620# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550#
+ m1_1540_1550# m1_1540_1550# m1_1540_1550# w_1650_2620# m2_n1840_n2910# m2_n1840_n2910#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# w_1650_2620# w_1650_2620# m2_n1840_n2910#
+ m1_1540_1550# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550#
+ m1_1540_1550# m1_1540_1550# m2_n1840_n2910# w_1686_386# m2_n1840_n2910# w_1650_2620#
+ w_1650_2620# w_1686_386# m2_n1840_n2910# m1_1540_1550# w_1650_2620# w_1650_2620#
+ m1_1540_1550# m2_n1840_n2910# m1_1540_1550# w_1686_386# m2_n1840_n2910# m1_1540_1550#
+ m1_1540_1550# m1_1540_1550# m2_n1840_n2910# w_1650_2620# w_1650_2620# m2_n1840_n2910#
+ w_1650_2620# m1_1540_1550# m1_1540_1550# m1_1540_1550# m1_1540_1550# m1_1540_1550#
+ m2_n1840_n2910# w_1650_2620# m1_1540_1550# m2_n1840_n2910# w_1686_386# w_1650_2620#
+ m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# m2_n1840_n2910# m1_1540_1550#
+ m1_1540_1550# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# w_1650_2620#
+ m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550# w_1650_2620# m1_1540_1550# w_1650_2620#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m2_n1840_n2910# w_1650_2620#
+ w_1686_386# w_1686_386# m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m1_1540_1550#
+ m1_1540_1550# m2_n1840_n2910# w_1650_2620# m1_1540_1550# w_1650_2620# m1_1540_1550#
+ w_1686_386# m2_n1840_n2910# w_1650_2620# m2_n1840_n2910# m1_1540_1550# m1_1540_1550#
+ m1_1540_1550# m2_n1840_n2910# w_1650_2620# m1_1540_1550# m1_1540_1550# m1_1540_1550#
+ w_1650_2620# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# m1_1540_1550# m1_1540_1550#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m1_1540_1550# w_1650_2620# m2_n1840_n2910#
+ m1_1540_1550# w_1650_2620# m1_1540_1550# m2_n1840_n2910# m2_n1840_n2910# m1_1540_1550#
+ m2_n1840_n2910# m1_1540_1550# m1_1540_1550# m2_n1840_n2910# w_1650_2620# m2_n1840_n2910#
+ m1_1540_1550# VSUBS m2_n1840_n2910# m1_1540_1550# m2_n1840_n2910# rf_transistors
Xsky130_fd_pr__cap_mim_m3_2_ZWVPUJ_0 m2_n1840_n2910# w_1650_2620# sky130_fd_pr__cap_mim_m3_2_ZWVPUJ
Xdis_tran_0 m2_n1840_n2910# m2_n1840_n2910# VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910#
+ m2_n1840_n2910# m2_n1840_n2910# m2_n1840_n2910# VSUBS VSUBS VSUBS m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# m2_n1840_n2910# VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910#
+ m2_n1840_n2910# m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# m1_n1960_n3240# m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910# VSUBS m1_n1960_n3240#
+ m2_n1840_n2910# VSUBS m2_n1840_n2910# VSUBS VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910#
+ VSUBS m2_n1840_n2910# m1_n1960_n3240# VSUBS VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910#
+ VSUBS m1_n1960_n3240# m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910#
+ m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910# m2_n1840_n2910# VSUBS VSUBS
+ VSUBS VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m2_n1840_n2910# m2_n1840_n2910#
+ VSUBS VSUBS m2_n1840_n2910# VSUBS m2_n1840_n2910# m1_n1960_n3240# VSUBS m2_n1840_n2910#
+ m2_n1840_n2910# VSUBS VSUBS VSUBS m2_n1840_n2910# VSUBS VSUBS m2_n1840_n2910# m2_n1840_n2910#
+ VSUBS dis_tran
Xfb_transistor_0 w_1686_386# w_1650_2620# m1_1850_2290# m2_1800_2380# w_1686_386#
+ m2_1800_2380# m1_1850_2290# m2_1800_2380# w_1686_386# w_1686_386# w_1650_2620# m2_1800_2380#
+ m2_1800_2380# w_1650_2620# w_1686_386# m1_1850_2290# m2_1800_2380# m1_1540_1550#
+ m2_1800_2380# w_1686_386# m2_1800_2380# m1_1850_2290# w_1686_386# m2_1800_2380#
+ w_1650_2620# m2_1800_2380# w_1686_386# m2_1800_2380# m2_1800_2380# w_1686_386# w_1686_386#
+ m2_1800_2380# w_1686_386# m2_1800_2380# m1_1850_2290# m1_1850_2290# m2_1800_2380#
+ w_1686_386# m2_1800_2380# m2_1800_2380# m1_1850_2290# w_1686_386# m2_1800_2380#
+ m2_1800_2380# w_1686_386# m1_1540_1550# m1_1850_2290# m2_1800_2380# m2_1800_2380#
+ w_1686_386# m1_1850_2290# w_1686_386# m1_1850_2290# w_1686_386# m2_1800_2380# w_1650_2620#
+ w_1650_2620# fb_transistor
.ends

.subckt sky130_fd_pr__pfet_01v8_GCYTE7 a_100_n50# w_n296_n269# a_n158_n50# a_n100_n147#
X0 a_100_n50# a_n100_n147# a_n158_n50# w_n296_n269# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_J5CT7Z c1_n1550_n1200# m3_n1650_n1300#
X0 c1_n1550_n1200# m3_n1650_n1300# sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=1.5e+07u
.ends

.subckt sky130_fd_pr__cap_var_lvt_MZUN4J a_n2040_n588# w_1507_n618# w_n2173_n618#
+ w_n333_n618# a_n1120_n588# w_587_n618# w_n1253_n618# a_n200_n588# a_1640_n588# a_720_n588#
X0 a_n200_n588# w_n333_n618# w_n333_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X1 a_n1120_n588# w_n1253_n618# w_n1253_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X2 a_720_n588# w_587_n618# w_587_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X3 a_1640_n588# w_1507_n618# w_1507_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
X4 a_n2040_n588# w_n2173_n618# w_n2173_n618# sky130_fd_pr__cap_var_lvt pd=2.194e+07u ps=0u ad=0p as=0p w=5e+06u l=2e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG#0 m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_SC2JGL a_15_n200# a_n177_n200# a_111_n200# a_159_n288#
+ a_63_222# a_n81_n200# a_n129_222# a_n269_n200# a_207_n200# a_n225_n288# a_n371_n374#
+ a_n33_n288#
X0 a_n81_n200# a_n129_222# a_n177_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_15_n200# a_n33_n288# a_n81_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X2 a_207_n200# a_159_n288# a_111_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n177_n200# a_n225_n288# a_n269_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X4 a_111_n200# a_63_222# a_15_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt tia_core VPP Out_2 Out_1 Disable_TIA I_Bias1 Out_ref VM39D Input VN
Xsky130_fd_pr__nfet_01v8_CDW43Z_0 VN Disable_TIA VN Disable_TIA_B sky130_fd_pr__nfet_01v8_CDW43Z
Xtia_cur_mirror_0 VN I_Bias1 VM6D I_Bias1 VN tia_cur_mirror
Xtia_one_tia_0 Disable_TIA_B VN Out_2 VM5D Input VPP I_Bias1 VM28D VN Out_1 tia_one_tia
Xtia_one_tia_1 Disable_TIA_B VN VM31D VM36D VM39D VPP I_Bias1 VM40D VN Out_ref tia_one_tia
Xsky130_fd_pr__pfet_01v8_GCYTE7_0 VPP VPP Disable_TIA_B Disable_TIA sky130_fd_pr__pfet_01v8_GCYTE7
Xsky130_fd_pr__cap_mim_m3_1_J5CT7Z_1 VN I_Bias1 sky130_fd_pr__cap_mim_m3_1_J5CT7Z
Xsky130_fd_pr__cap_mim_m3_1_J5CT7Z_0 VN I_Bias1 sky130_fd_pr__cap_mim_m3_1_J5CT7Z
Xsky130_fd_pr__cap_var_lvt_MZUN4J_0 Disable_TIA_B VN VN VN Disable_TIA_B VN VN Disable_TIA_B
+ Disable_TIA_B Disable_TIA_B sky130_fd_pr__cap_var_lvt_MZUN4J
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_0 VN VPP sky130_fd_pr__cap_mim_m3_2_LJ5JLG#0
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_1 VN VPP sky130_fd_pr__cap_mim_m3_2_LJ5JLG#0
Xsky130_fd_pr__nfet_01v8_SC2JGL_0 VN VN I_Bias1 Disable_TIA Disable_TIA I_Bias1 Disable_TIA
+ I_Bias1 VN Disable_TIA VN Disable_TIA sky130_fd_pr__nfet_01v8_SC2JGL
.ends

.subckt sky130_fd_pr__nfet_01v8_HR8DH9 a_262_n288# a_n328_n288# a_n501_n200# a_616_n288#
+ a_561_n200# a_144_n288# a_n839_n374# a_n383_n200# a_498_n288# a_n737_n200# a_443_n200#
+ a_n265_n200# a_n619_n200# a_26_n288# a_325_n200# a_n682_n288# a_679_n200# a_n147_n200#
+ a_207_n200# a_n210_n288# a_n564_n288# a_n29_n200# a_380_n288# a_n92_n288# a_89_n200#
+ a_n446_n288#
X0 a_n29_n200# a_n92_n288# a_n147_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X1 a_n619_n200# a_n682_n288# a_n737_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X2 a_325_n200# a_262_n288# a_207_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X3 a_561_n200# a_498_n288# a_443_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X4 a_n265_n200# a_n328_n288# a_n383_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X5 a_89_n200# a_26_n288# a_n29_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X6 a_207_n200# a_144_n288# a_89_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X7 a_n501_n200# a_n564_n288# a_n619_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X8 a_n147_n200# a_n210_n288# a_n265_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X9 a_679_n200# a_616_n288# a_561_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X10 a_443_n200# a_380_n288# a_325_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X11 a_n383_n200# a_n446_n288# a_n501_n200# a_n839_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
.ends

.subckt sky130_fd_pr__nfet_01v8_XZXALN a_n129_727# a_n129_109# a_n369_21# a_n177_n1215#
+ a_n605_n1127# a_n465_n597# a_255_n509# a_n561_n1215# a_n707_n1301# a_495_n705# a_n273_639#
+ a_15_1149# a_399_21# a_n561_1149# a_447_727# a_n81_531# a_447_109# a_399_n1215#
+ a_n177_1149# a_351_n509# a_n417_n509# a_n177_n87# a_n321_727# a_n321_109# a_111_n597#
+ a_63_n1127# a_n273_531# a_n273_n597# a_n513_n509# a_n33_n1127# a_n129_n509# a_159_727#
+ a_159_109# a_303_n705# a_63_n509# a_n417_n1127# a_n129_n1127# a_n465_639# a_n513_n1127#
+ a_n225_n1127# a_n321_n1127# a_n369_n87# a_n225_n509# a_n465_n705# a_n513_727# a_n513_109#
+ a_n465_531# a_159_n1127# a_447_n1127# a_255_n1127# a_543_n1127# a_351_n1127# a_351_727#
+ a_351_109# a_n321_n509# a_n33_727# a_n33_109# a_399_1149# a_n81_n597# a_111_n705#
+ a_n561_n87# a_n225_727# a_n225_109# a_495_639# a_n273_n705# a_15_n1215# a_111_639#
+ a_n561_21# a_n177_21# a_n33_n509# a_495_n597# a_207_21# a_399_n87# a_543_727# a_543_109#
+ a_495_531# a_111_531# a_n605_n509# a_63_727# a_63_109# a_447_n509# a_15_n87# a_207_1149#
+ a_n605_727# a_15_21# a_n605_109# a_n417_727# a_n417_109# a_303_639# a_207_n1215#
+ a_n369_1149# a_255_727# a_255_109# a_543_n509# a_159_n509# a_n81_n705# a_207_n87#
+ a_303_n597# a_303_531# a_n81_639# a_n369_n1215#
X0 a_n129_n509# a_n177_n87# a_n225_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n321_n1127# a_n369_n1215# a_n417_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_n417_n509# a_n465_n597# a_n513_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n33_727# a_n81_639# a_n129_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_351_727# a_303_639# a_255_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_159_727# a_111_639# a_63_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_255_727# a_207_1149# a_159_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 a_447_727# a_399_1149# a_351_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X8 a_543_727# a_495_639# a_447_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X9 a_63_n1127# a_15_n1215# a_n33_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_159_n1127# a_111_n705# a_63_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_n33_109# a_n81_531# a_n129_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_n33_n509# a_n81_n597# a_n129_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X13 a_351_n509# a_303_n597# a_255_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X14 a_n321_727# a_n369_1149# a_n417_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X15 a_255_n1127# a_207_n1215# a_159_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X16 a_n513_727# a_n561_1149# a_n605_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X17 a_n417_727# a_n465_639# a_n513_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 a_n225_727# a_n273_639# a_n321_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X19 a_n129_727# a_n177_1149# a_n225_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 a_255_109# a_207_21# a_159_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X21 a_351_109# a_303_531# a_255_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X22 a_543_109# a_495_531# a_447_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X23 a_n417_n1127# a_n465_n705# a_n513_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X24 a_159_109# a_111_531# a_63_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X25 a_447_109# a_399_21# a_351_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 a_n513_n1127# a_n561_n1215# a_n605_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X27 a_351_n1127# a_303_n705# a_255_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X28 a_n513_109# a_n561_21# a_n605_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X29 a_n321_109# a_n369_21# a_n417_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X30 a_n225_109# a_n273_531# a_n321_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X31 a_n417_109# a_n465_531# a_n513_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 a_n129_109# a_n177_21# a_n225_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 a_255_n509# a_207_n87# a_159_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X34 a_n321_n509# a_n369_n87# a_n417_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X35 a_63_727# a_15_1149# a_n33_727# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 a_543_n509# a_495_n597# a_447_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X37 a_n33_n1127# a_n81_n705# a_n129_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X38 a_63_109# a_15_21# a_n33_109# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X39 a_159_n509# a_111_n597# a_63_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X40 a_n225_n509# a_n273_n597# a_n321_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X41 a_447_n509# a_399_n87# a_351_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X42 a_n129_n1127# a_n177_n1215# a_n225_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X43 a_447_n1127# a_399_n1215# a_351_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X44 a_n513_n509# a_n561_n87# a_n605_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X45 a_63_n509# a_15_n87# a_n33_n509# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 a_n225_n1127# a_n273_n705# a_n321_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 a_543_n1127# a_495_n705# a_447_n1127# a_n707_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt lvds_currm_n m1_76_644# m1_n20_420# a_42_42# VSUBS
Xsky130_fd_pr__nfet_01v8_HR8DH9_0 a_42_42# a_42_42# VSUBS a_42_42# m1_n20_420# a_42_42#
+ VSUBS m1_n20_420# a_42_42# VSUBS VSUBS VSUBS m1_n20_420# a_42_42# m1_n20_420# a_42_42#
+ VSUBS m1_n20_420# VSUBS a_42_42# a_42_42# VSUBS a_42_42# a_42_42# m1_n20_420# a_42_42#
+ sky130_fd_pr__nfet_01v8_HR8DH9
Xsky130_fd_pr__nfet_01v8_XZXALN_0 m1_76_644# m1_76_644# a_42_42# a_42_42# m1_n20_420#
+ a_42_42# m1_76_644# a_42_42# VSUBS a_42_42# a_42_42# a_42_42# a_42_42# a_42_42#
+ m1_76_644# a_42_42# m1_76_644# a_42_42# a_42_42# m1_n20_420# m1_n20_420# a_42_42#
+ m1_76_644# m1_76_644# a_42_42# m1_76_644# a_42_42# a_42_42# m1_76_644# m1_n20_420#
+ m1_76_644# m1_n20_420# m1_n20_420# a_42_42# m1_76_644# m1_n20_420# m1_76_644# a_42_42#
+ m1_76_644# m1_n20_420# m1_76_644# a_42_42# m1_n20_420# a_42_42# m1_76_644# m1_76_644#
+ a_42_42# m1_n20_420# m1_76_644# m1_76_644# m1_n20_420# m1_n20_420# m1_n20_420# m1_n20_420#
+ m1_76_644# m1_n20_420# m1_n20_420# a_42_42# a_42_42# a_42_42# a_42_42# m1_n20_420#
+ m1_n20_420# a_42_42# a_42_42# a_42_42# a_42_42# a_42_42# a_42_42# m1_n20_420# a_42_42#
+ a_42_42# a_42_42# m1_n20_420# m1_n20_420# a_42_42# a_42_42# m1_n20_420# m1_76_644#
+ m1_76_644# m1_76_644# a_42_42# a_42_42# m1_n20_420# a_42_42# m1_n20_420# m1_n20_420#
+ m1_n20_420# a_42_42# a_42_42# a_42_42# m1_76_644# m1_76_644# m1_n20_420# m1_n20_420#
+ a_42_42# a_42_42# a_42_42# a_42_42# a_42_42# a_42_42# sky130_fd_pr__nfet_01v8_XZXALN
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL a_n194_n1432# a_n324_n1562# a_n194_1000#
+ a_124_n1432# a_124_1000#
X0 a_124_n1432# a_124_1000# a_n324_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
X1 a_n194_n1432# a_n194_1000# a_n324_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
.ends

.subckt sky130_fd_sc_hs__inv_16 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=2.7216e+12p pd=2.278e+07u as=3.4272e+12p ps=2.628e+07u w=1.12e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=1.6576e+12p pd=1.632e+07u as=2.2718e+12p ps=1.946e+07u w=740000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X27 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X30 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_RS2YEK a_283_1000# a_n353_n1432# a_n35_n1432#
+ a_n35_1000# a_n483_n1562# a_n353_1000# a_283_n1432#
X0 a_n353_n1432# a_n353_1000# a_n483_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
X1 a_283_n1432# a_283_1000# a_n483_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
X2 a_n35_n1432# a_n35_1000# a_n483_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_8DK6RJ a_n321_n518# a_255_n1154# a_543_n1154# a_n369_21#
+ a_n33_118# a_351_754# a_351_n1154# a_n81_657# a_n33_754# a_495_n723# a_n369_n1251#
+ a_n177_n1251# a_n561_n1251# a_399_21# a_n225_118# w_n743_n1373# a_n273_657# a_n225_754#
+ a_n177_n87# a_15_1185# a_n33_n518# a_n561_1185# a_303_n615# a_n177_1185# a_399_n1251#
+ a_n465_549# a_543_118# a_543_754# a_n465_n615# a_n605_n518# a_63_118# a_447_n518#
+ a_63_754# a_n605_118# a_n417_118# a_303_n723# a_n465_657# a_n605_754# a_n417_754#
+ a_n369_n87# a_255_118# a_543_n518# a_159_n518# a_n465_n723# a_111_n615# a_255_754#
+ a_495_549# a_111_549# a_n273_n615# a_n129_118# a_255_n518# a_n129_754# a_n561_n87#
+ a_n605_n1154# a_111_n723# a_399_1185# a_n561_21# a_447_118# a_n177_21# a_495_657#
+ a_351_n518# a_n417_n518# a_111_657# a_447_754# a_n273_n723# a_207_21# a_399_n87#
+ a_15_n1251# a_n321_118# a_n321_754# a_303_549# a_63_n1154# a_n513_n518# a_n129_n518#
+ a_n81_n615# a_15_n87# a_15_21# a_n33_n1154# a_159_118# a_63_n518# a_159_754# a_207_1185#
+ a_n417_n1154# a_n129_n1154# a_n513_n1154# a_n225_n1154# a_n81_549# a_303_657# a_n321_n1154#
+ a_n225_n518# a_495_n615# a_n513_118# a_207_n87# a_n81_n723# a_n513_754# a_207_n1251#
+ a_n369_1185# a_n273_549# a_159_n1154# a_447_n1154# a_351_118#
X0 a_447_n518# a_399_n87# a_351_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n513_n518# a_n561_n87# a_n605_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X2 a_63_n518# a_15_n87# a_n33_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n33_754# a_n81_657# a_n129_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_351_754# a_303_657# a_255_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_159_754# a_111_657# a_63_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_255_754# a_207_1185# a_159_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 a_447_754# a_399_1185# a_351_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X8 a_543_754# a_495_657# a_447_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X9 a_63_n1154# a_15_n1251# a_n33_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_159_n1154# a_111_n723# a_63_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_n129_n518# a_n177_n87# a_n225_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_n513_754# a_n561_1185# a_n605_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X13 a_n321_754# a_n369_1185# a_n417_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X14 a_n225_754# a_n273_657# a_n321_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X15 a_255_n1154# a_207_n1251# a_159_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X16 a_n417_754# a_n465_657# a_n513_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 a_n129_754# a_n177_1185# a_n225_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 a_n417_n518# a_n465_n615# a_n513_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X19 a_n417_n1154# a_n465_n723# a_n513_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X20 a_351_n1154# a_303_n723# a_255_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X21 a_n513_n1154# a_n561_n1251# a_n605_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X22 a_63_754# a_15_1185# a_n33_754# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 a_n33_n518# a_n81_n615# a_n129_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 a_351_n518# a_303_n615# a_255_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X25 a_n33_118# a_n81_549# a_n129_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X26 a_351_118# a_303_549# a_255_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X27 a_159_118# a_111_549# a_63_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X28 a_255_118# a_207_21# a_159_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 a_447_118# a_399_21# a_351_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X30 a_543_118# a_495_549# a_447_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X31 a_n33_n1154# a_n81_n723# a_n129_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X32 a_n513_118# a_n561_21# a_n605_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X33 a_n321_118# a_n369_21# a_n417_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X34 a_n225_118# a_n273_549# a_n321_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X35 a_n417_118# a_n465_549# a_n513_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 a_n129_118# a_n177_21# a_n225_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 a_255_n518# a_207_n87# a_159_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X38 a_n129_n1154# a_n177_n1251# a_n225_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X39 a_447_n1154# a_399_n1251# a_351_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X40 a_n321_n518# a_n369_n87# a_n417_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X41 a_543_n518# a_495_n615# a_447_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X42 a_n225_n1154# a_n273_n723# a_n321_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X43 a_543_n1154# a_495_n723# a_447_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X44 a_n321_n1154# a_n369_n1251# a_n417_n1154# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X45 a_63_118# a_15_21# a_n33_118# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 a_159_n518# a_111_n615# a_63_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 a_n225_n518# a_n273_n615# a_n321_n518# w_n743_n1373# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_9Z5L4S a_n383_n518# a_498_n615# a_380_21# a_n92_21#
+ a_n737_n518# a_325_118# a_443_n518# a_n265_n518# a_89_118# a_n619_n518# a_26_n615#
+ a_n265_118# a_n501_118# a_679_n518# a_325_n518# a_n682_n615# a_n147_n518# a_443_118#
+ a_26_21# a_207_n518# a_n210_n615# a_n564_n615# a_n328_21# a_n383_118# a_n446_21#
+ a_n29_n518# a_n564_21# a_n619_118# a_n682_21# a_380_n615# a_n92_n615# a_89_n518#
+ a_n446_n615# a_561_118# a_n210_21# a_262_n615# a_n328_n615# a_n29_118# a_616_21#
+ a_498_21# a_207_118# a_n737_118# a_n501_n518# a_616_n615# w_n875_n737# a_144_21#
+ a_561_n518# a_144_n615# a_679_118# a_n147_118# a_262_21#
X0 a_n383_118# a_n446_21# a_n501_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X1 a_679_n518# a_616_n615# a_561_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X2 a_n29_118# a_n92_21# a_n147_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X3 a_n265_118# a_n328_21# a_n383_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X4 a_443_n518# a_380_n615# a_325_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X5 a_89_118# a_26_21# a_n29_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X6 a_n383_n518# a_n446_n615# a_n501_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X7 a_n147_118# a_n210_21# a_n265_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X8 a_679_118# a_616_21# a_561_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X9 a_443_118# a_380_21# a_325_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X10 a_n619_n518# a_n682_n615# a_n737_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X11 a_n29_n518# a_n92_n615# a_n147_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X12 a_561_118# a_498_21# a_443_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X13 a_325_n518# a_262_n615# a_207_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X14 a_325_118# a_262_21# a_207_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X15 a_561_n518# a_498_n615# a_443_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X16 a_n265_n518# a_n328_n615# a_n383_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X17 a_n619_118# a_n682_21# a_n737_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X18 a_207_118# a_144_21# a_89_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 a_n501_118# a_n564_21# a_n619_118# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X20 a_89_n518# a_26_n615# a_n29_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X21 a_207_n518# a_144_n615# a_89_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X22 a_n501_n518# a_n564_n615# a_n619_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X23 a_n147_n518# a_n210_n615# a_n265_n518# w_n875_n737# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
.ends

.subckt lvds_currm_p a_112_112# m1_60_208# m1_60_1070# w_112_640#
Xsky130_fd_pr__pfet_01v8_8DK6RJ_0 m1_60_208# m1_60_1070# m1_60_208# a_112_112# m1_60_1070#
+ m1_60_1070# m1_60_208# a_112_112# m1_60_1070# a_112_112# a_112_112# a_112_112# a_112_112#
+ a_112_112# m1_60_1070# w_112_640# a_112_112# m1_60_1070# a_112_112# a_112_112# m1_60_1070#
+ a_112_112# a_112_112# a_112_112# a_112_112# a_112_112# m1_60_1070# m1_60_1070# a_112_112#
+ m1_60_1070# m1_60_208# m1_60_208# m1_60_208# m1_60_1070# m1_60_1070# a_112_112#
+ a_112_112# m1_60_1070# m1_60_1070# a_112_112# m1_60_208# m1_60_1070# m1_60_1070#
+ a_112_112# a_112_112# m1_60_208# a_112_112# a_112_112# a_112_112# m1_60_208# m1_60_208#
+ m1_60_208# a_112_112# m1_60_208# a_112_112# a_112_112# a_112_112# m1_60_208# a_112_112#
+ a_112_112# m1_60_1070# m1_60_1070# a_112_112# m1_60_208# a_112_112# a_112_112# a_112_112#
+ a_112_112# m1_60_208# m1_60_208# a_112_112# m1_60_1070# m1_60_208# m1_60_208# a_112_112#
+ a_112_112# a_112_112# m1_60_208# m1_60_1070# m1_60_208# m1_60_1070# a_112_112# m1_60_208#
+ m1_60_1070# m1_60_1070# m1_60_208# a_112_112# a_112_112# m1_60_1070# m1_60_1070#
+ a_112_112# m1_60_208# a_112_112# a_112_112# m1_60_208# a_112_112# a_112_112# a_112_112#
+ m1_60_208# m1_60_1070# m1_60_1070# sky130_fd_pr__pfet_01v8_8DK6RJ
Xsky130_fd_pr__pfet_01v8_9Z5L4S_0 w_112_640# a_112_112# a_112_112# a_112_112# m1_60_1070#
+ w_112_640# m1_60_1070# m1_60_1070# w_112_640# w_112_640# a_112_112# m1_60_1070#
+ m1_60_1070# m1_60_1070# w_112_640# a_112_112# w_112_640# m1_60_1070# a_112_112#
+ m1_60_1070# a_112_112# a_112_112# a_112_112# w_112_640# a_112_112# m1_60_1070# a_112_112#
+ w_112_640# a_112_112# a_112_112# a_112_112# w_112_640# a_112_112# w_112_640# a_112_112#
+ a_112_112# a_112_112# m1_60_1070# a_112_112# a_112_112# m1_60_1070# m1_60_1070#
+ m1_60_1070# a_112_112# w_112_640# a_112_112# w_112_640# a_112_112# m1_60_1070# w_112_640#
+ a_112_112# sky130_fd_pr__pfet_01v8_9Z5L4S
.ends

.subckt sky130_fd_pr__pfet_01v8_VCB4SW a_351_436# a_n81_339# a_n513_n200# a_n321_n836#
+ a_n1329_n297# a_n753_867# a_n33_436# a_n129_n200# a_n945_n405# a_n657_n933# a_831_436#
+ a_15_867# a_639_n836# a_1311_436# a_63_n200# a_1215_n200# a_1023_n836# a_n1041_231#
+ a_879_339# a_n1281_n836# a_1167_n297# a_n1089_n200# a_591_867# a_n273_339# a_n225_436#
+ a_15_n297# a_n81_231# a_n225_n200# a_n1089_436# a_n561_n297# a_591_n405# a_n177_n297#
+ a_n705_436# a_207_867# a_927_n200# a_1311_n200# a_n33_n836# a_735_n836# a_n1233_339#
+ a_303_n933# a_879_231# a_n1185_n200# a_207_n405# a_1359_n405# a_n273_231# a_543_436#
+ a_n1469_n836# a_1071_339# a_n945_867# a_1023_436# a_n321_n200# a_n897_n836# a_n1137_n297#
+ a_n753_n405# a_n465_n933# a_n369_n405# a_831_n836# a_n1233_231# a_63_436# a_975_n297#
+ a_639_n200# a_1023_n200# a_447_n836# a_783_867# a_n1281_n200# a_n1281_436# a_n465_339#
+ a_n417_436# a_1071_231# a_n1469_436# a_n993_n836# a_n1425_n933# a_n1329_n405# a_n177_867#
+ a_n1425_339# a_255_436# a_n33_n200# a_735_n200# a_543_n836# a_n609_n836# a_159_n836#
+ a_111_n933# a_879_n933# a_1263_n933# a_n465_231# a_1167_n405# a_735_436# a_1263_339#
+ a_n1469_n200# a_n1137_867# a_1215_436# a_n897_n200# a_15_n405# a_n993_436# a_n561_n405#
+ a_n273_n933# a_n177_n405# a_n1425_231# a_831_n200# a_n129_436# a_n705_n836# a_975_867#
+ a_783_n297# a_447_n200# a_255_n836# a_399_n297# a_n657_339# a_n609_436# a_1263_231#
+ a_1407_n836# a_n993_n200# a_n1233_n933# a_n369_867# a_n1137_n405# a_495_339# a_447_436#
+ a_111_339# a_543_n200# a_n801_n836# a_351_n836# a_n609_n200# a_n417_n836# a_159_n200#
+ a_975_n405# a_n945_n297# a_n657_231# a_687_n933# a_927_436# a_1071_n933# a_n1329_867#
+ a_1407_436# a_n321_436# a_1119_n836# a_n1377_n836# a_n1185_436# a_495_231# a_n801_436#
+ a_1167_867# a_111_231# a_n849_339# a_n705_n200# a_255_n200# a_n513_n836# a_n129_n836#
+ a_591_n297# a_n81_n933# a_n561_867# a_n849_n933# a_1407_n200# a_1215_n836# a_159_436#
+ a_63_n836# a_207_n297# a_1359_n297# w_n1607_n1055# a_n1089_n836# a_687_339# a_n1041_n933#
+ a_639_436# a_303_339# a_n801_n200# a_1119_436# a_351_n200# a_n849_231# a_n417_n200#
+ a_n225_n836# a_n753_n297# a_783_n405# a_n897_436# a_399_867# a_495_n933# a_n369_n297#
+ a_399_n405# a_n513_436# a_927_n836# a_1311_n836# a_1119_n200# a_n1377_436# a_n1041_339#
+ a_n1377_n200# a_n1185_n836# a_687_231# a_1359_867# a_303_231#
X0 a_n1281_n200# a_n1329_n297# a_n1377_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n609_n200# a_n657_231# a_n705_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_n417_n836# a_n465_n933# a_n513_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_927_n200# a_879_231# a_831_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_639_n836# a_591_n405# a_543_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_927_436# a_879_339# a_831_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_1023_436# a_975_867# a_927_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X7 a_n897_n200# a_n945_n297# a_n993_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X8 a_n705_n836# a_n753_n405# a_n801_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X9 a_255_n200# a_207_n297# a_159_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_1215_n200# a_1167_n297# a_1119_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X11 a_1119_436# a_1071_339# a_1023_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X12 a_1215_436# a_1167_867# a_1119_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X13 a_1311_436# a_1263_339# a_1215_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X14 a_1407_436# a_1359_867# a_1311_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X15 a_n321_n200# a_n369_n297# a_n417_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X16 a_1023_n836# a_975_n405# a_927_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17 a_n1185_n200# a_n1233_231# a_n1281_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X18 a_543_n200# a_495_231# a_447_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X19 a_1311_n836# a_1263_n933# a_1215_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X20 a_n993_n836# a_n1041_n933# a_n1089_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X21 a_n33_n836# a_n81_n933# a_n129_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X22 a_351_n836# a_303_n933# a_255_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X23 a_n33_436# a_n81_339# a_n129_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X24 a_351_436# a_303_339# a_255_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X25 a_831_n200# a_783_n297# a_735_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X26 a_159_436# a_111_339# a_63_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X27 a_255_436# a_207_867# a_159_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 a_447_436# a_399_867# a_351_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X29 a_543_436# a_495_339# a_447_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X30 a_639_436# a_591_867# a_543_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X31 a_735_436# a_687_339# a_639_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X32 a_831_436# a_783_867# a_735_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 a_159_n200# a_111_231# a_63_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X34 a_1119_n200# a_1071_231# a_1023_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X35 a_n1281_n836# a_n1329_n405# a_n1377_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X36 a_n609_n836# a_n657_n933# a_n705_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X37 a_n1377_436# a_n1425_339# a_n1469_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X38 a_n1281_436# a_n1329_867# a_n1377_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X39 a_n1185_436# a_n1233_339# a_n1281_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X40 a_n1089_436# a_n1137_867# a_n1185_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X41 a_n993_436# a_n1041_339# a_n1089_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X42 a_n225_n200# a_n273_231# a_n321_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X43 a_n897_n836# a_n945_n405# a_n993_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X44 a_927_n836# a_879_n933# a_831_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X45 a_n801_436# a_n849_339# a_n897_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X46 a_n513_436# a_n561_867# a_n609_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X47 a_n321_436# a_n369_867# a_n417_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X48 a_n225_436# a_n273_339# a_n321_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X49 a_n1089_n200# a_n1137_n297# a_n1185_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X50 a_447_n200# a_399_n297# a_351_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X51 a_1407_n200# a_1359_n297# a_1311_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X52 a_1215_n836# a_1167_n405# a_1119_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X53 a_n897_436# a_n945_867# a_n993_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 a_n705_436# a_n753_867# a_n801_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X55 a_n609_436# a_n657_339# a_n705_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X56 a_n417_436# a_n465_339# a_n513_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X57 a_n129_436# a_n177_867# a_n225_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X58 a_255_n836# a_207_n405# a_159_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X59 a_n513_n200# a_n561_n297# a_n609_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X60 a_63_n200# a_15_n297# a_n33_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X61 a_n321_n836# a_n369_n405# a_n417_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X62 a_n1377_n200# a_n1425_231# a_n1469_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X63 a_735_n200# a_687_231# a_639_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X64 a_543_n836# a_495_n933# a_447_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X65 a_n801_n200# a_n849_231# a_n897_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X66 a_n1185_n836# a_n1233_n933# a_n1281_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X67 a_n129_n200# a_n177_n297# a_n225_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X68 a_831_n836# a_783_n405# a_735_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X69 a_1119_n836# a_1071_n933# a_1023_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X70 a_63_436# a_15_867# a_n33_436# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 a_159_n836# a_111_n933# a_63_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X72 a_n417_n200# a_n465_231# a_n513_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X73 a_n225_n836# a_n273_n933# a_n321_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X74 a_639_n200# a_591_n297# a_543_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X75 a_447_n836# a_399_n405# a_351_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X76 a_1407_n836# a_1359_n405# a_1311_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X77 a_n705_n200# a_n753_n297# a_n801_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 a_n1089_n836# a_n1137_n405# a_n1185_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 a_n513_n836# a_n561_n405# a_n609_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X80 a_63_n836# a_15_n405# a_n33_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 a_1023_n200# a_975_n297# a_927_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 a_n1377_n836# a_n1425_n933# a_n1469_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X83 a_735_n836# a_687_n933# a_639_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 a_n801_n836# a_n849_n933# a_n897_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X85 a_351_n200# a_303_231# a_255_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 a_1311_n200# a_1263_231# a_1215_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 a_n993_n200# a_n1041_231# a_n1089_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X88 a_n33_n200# a_n81_231# a_n129_n200# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 a_n129_n836# a_n177_n405# a_n225_n836# w_n1607_n1055# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt lvds_switch_p m1_178_212# m1_274_438# m1_178_1074# m1_274_848# m1_178_1484#
+ a_230_644# m1_274_1710# w_230_752#
Xsky130_fd_pr__pfet_01v8_VCB4SW_0 m1_274_1710# a_230_644# m1_178_1074# m1_178_212#
+ a_230_644# a_230_644# m1_274_1710# m1_178_1074# a_230_644# a_230_644# m1_178_1484#
+ a_230_644# m1_178_212# m1_274_1710# m1_178_1074# m1_178_1074# m1_178_212# a_230_644#
+ a_230_644# m1_178_212# a_230_644# m1_178_1074# a_230_644# a_230_644# m1_274_1710#
+ a_230_644# a_230_644# m1_274_848# m1_178_1484# a_230_644# a_230_644# a_230_644#
+ m1_178_1484# a_230_644# m1_274_848# m1_274_848# m1_274_438# m1_274_438# a_230_644#
+ a_230_644# a_230_644# m1_274_848# a_230_644# a_230_644# a_230_644# m1_274_1710#
+ m1_178_212# a_230_644# a_230_644# m1_178_1484# m1_178_1074# m1_178_212# a_230_644#
+ a_230_644# a_230_644# a_230_644# m1_178_212# a_230_644# m1_178_1484# a_230_644#
+ m1_178_1074# m1_178_1074# m1_178_212# a_230_644# m1_178_1074# m1_178_1484# a_230_644#
+ m1_274_1710# a_230_644# m1_178_1484# m1_274_438# a_230_644# a_230_644# a_230_644#
+ a_230_644# m1_178_1484# m1_274_848# m1_274_848# m1_274_438# m1_274_438# m1_274_438#
+ a_230_644# a_230_644# a_230_644# a_230_644# a_230_644# m1_274_1710# a_230_644# m1_178_1074#
+ a_230_644# m1_178_1484# m1_178_1074# a_230_644# m1_274_1710# a_230_644# a_230_644#
+ a_230_644# a_230_644# m1_178_1074# m1_178_1484# m1_178_212# a_230_644# a_230_644#
+ m1_178_1074# m1_178_212# a_230_644# a_230_644# m1_274_1710# a_230_644# m1_178_212#
+ m1_274_848# a_230_644# a_230_644# a_230_644# a_230_644# m1_178_1484# a_230_644#
+ m1_274_848# m1_274_438# m1_274_438# m1_274_848# m1_274_438# m1_274_848# a_230_644#
+ a_230_644# a_230_644# a_230_644# m1_274_1710# a_230_644# a_230_644# m1_178_1484#
+ m1_178_1484# m1_274_438# m1_274_438# m1_274_1710# a_230_644# m1_274_1710# a_230_644#
+ a_230_644# a_230_644# m1_178_1074# m1_178_1074# m1_178_212# m1_178_212# a_230_644#
+ a_230_644# a_230_644# a_230_644# m1_178_1074# m1_178_212# m1_274_1710# m1_178_212#
+ a_230_644# a_230_644# w_230_752# m1_178_212# a_230_644# a_230_644# m1_178_1484#
+ a_230_644# m1_274_848# m1_274_1710# m1_274_848# a_230_644# m1_274_848# m1_274_438#
+ a_230_644# a_230_644# m1_178_1484# a_230_644# a_230_644# a_230_644# a_230_644# m1_178_1484#
+ m1_274_438# m1_274_438# m1_274_848# m1_274_1710# a_230_644# m1_274_848# m1_274_438#
+ a_230_644# a_230_644# a_230_644# sky130_fd_pr__pfet_01v8_VCB4SW
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_N3PKNJ c1_n3050_n1000# m3_n3150_n1100#
X0 c1_n3050_n1000# m3_n3150_n1100# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_RE4MKQ a_n1041_109# a_n993_531# a_1119_n597# a_n1229_109#
+ a_n753_n509# a_n81_109# a_n369_n509# a_n705_21# a_399_109# a_303_n509# a_831_n87#
+ a_n609_531# a_879_109# a_n273_109# a_n465_n509# a_n753_109# a_n1089_n87# a_927_531#
+ a_15_109# a_n705_n87# a_n1089_21# a_n225_n597# a_1167_n509# a_927_n597# a_n1185_531#
+ a_591_109# a_15_n509# a_n801_531# a_n1185_n597# a_1071_109# a_n561_n509# a_n177_n509#
+ a_1023_n87# a_n321_21# a_207_109# a_111_n509# a_879_n509# a_159_531# a_639_21# a_63_n87#
+ a_n465_109# a_n1137_n509# a_n273_n509# a_1119_531# a_n945_109# a_975_n509# a_255_n87#
+ a_783_109# a_n33_n597# a_735_n597# a_n897_21# a_351_531# a_n1331_n683# a_n33_531#
+ a_n177_109# a_687_n509# a_1071_n509# a_n129_n87# a_255_21# a_n657_109# a_n225_531#
+ a_n1137_109# a_495_109# a_111_109# a_n993_n597# a_n81_n509# a_783_n509# a_n513_21#
+ a_447_n87# a_n849_n509# a_399_n509# a_n129_21# a_1023_21# a_975_109# a_63_21# a_543_n597#
+ a_n609_n597# a_159_n597# a_543_531# a_n1041_n509# a_n321_n87# a_n369_109# a_n945_n509#
+ a_495_n509# a_n849_109# a_n417_531# a_687_109# a_n1229_n509# a_303_109# a_1167_109#
+ a_639_n87# a_591_n509# a_n657_n509# a_n561_109# a_831_21# a_n897_n87# a_n801_n597#
+ a_351_n597# a_447_21# a_735_531# a_n417_n597# a_207_n509# a_n513_n87#
X0 a_399_n509# a_351_n597# a_303_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n81_109# a_n129_21# a_n177_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_111_109# a_63_21# a_15_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n465_n509# a_n513_n87# a_n561_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n273_109# a_n321_21# a_n369_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_n177_109# a_n225_531# a_n273_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 a_687_n509# a_639_n87# a_591_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_n753_n509# a_n801_n597# a_n849_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X8 a_975_n509# a_927_n597# a_879_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X9 a_n81_n509# a_n129_n87# a_n177_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_15_n509# a_n33_n597# a_n81_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_n1041_n509# a_n1089_n87# a_n1137_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_n369_n509# a_n417_n597# a_n465_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X13 a_n657_n509# a_n705_n87# a_n753_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X14 a_879_n509# a_831_n87# a_783_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X15 a_n945_n509# a_n993_n597# a_n1041_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X16 a_1167_n509# a_1119_n597# a_1071_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17 a_303_n509# a_255_n87# a_207_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X18 a_n273_n509# a_n321_n87# a_n369_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X19 a_591_n509# a_543_n597# a_495_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X20 a_n849_n509# a_n897_n87# a_n945_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 a_303_109# a_255_21# a_207_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X22 a_591_109# a_543_531# a_495_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X23 a_207_109# a_159_531# a_111_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 a_399_109# a_351_531# a_303_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X25 a_495_109# a_447_21# a_399_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 a_687_109# a_639_21# a_591_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X27 a_783_109# a_735_531# a_687_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X28 a_975_109# a_927_531# a_879_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X29 a_n177_n509# a_n225_n597# a_n273_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 a_207_n509# a_159_n597# a_111_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X31 a_n1041_109# a_n1089_21# a_n1137_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X32 a_879_109# a_831_21# a_783_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 a_n1137_109# a_n1185_531# a_n1229_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X34 a_n1137_n509# a_n1185_n597# a_n1229_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X35 a_495_n509# a_447_n87# a_399_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 a_n561_109# a_n609_531# a_n657_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X37 a_1071_109# a_1023_21# a_975_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X38 a_n945_109# a_n993_531# a_n1041_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X39 a_n753_109# a_n801_531# a_n849_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X40 a_n657_109# a_n705_21# a_n753_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X41 a_n465_109# a_n513_21# a_n561_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X42 a_n369_109# a_n417_531# a_n465_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X43 a_1167_109# a_1119_531# a_1071_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X44 a_n561_n509# a_n609_n597# a_n657_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X45 a_111_n509# a_63_n87# a_15_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 a_n849_109# a_n897_21# a_n945_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 a_783_n509# a_735_n597# a_687_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X48 a_15_109# a_n33_531# a_n81_109# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 a_1071_n509# a_1023_n87# a_975_n509# a_n1331_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt lvds_nswitch m1_30_728# m1_126_952# m1_30_110# a_82_22# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_RE4MKQ_0 m1_30_728# a_82_22# a_82_22# m1_30_728# m1_30_728#
+ m1_30_728# m1_30_728# a_82_22# m1_126_952# m1_30_110# a_82_22# a_82_22# m1_30_728#
+ m1_30_728# m1_30_110# m1_126_952# a_82_22# a_82_22# m1_126_952# a_82_22# a_82_22#
+ a_82_22# m1_30_728# a_82_22# a_82_22# m1_126_952# m1_30_728# a_82_22# a_82_22# m1_30_728#
+ m1_30_728# m1_30_728# a_82_22# a_82_22# m1_126_952# m1_30_110# m1_30_110# a_82_22#
+ a_82_22# a_82_22# m1_30_728# m1_30_728# m1_30_110# a_82_22# m1_126_952# m1_30_728#
+ a_82_22# m1_126_952# a_82_22# a_82_22# a_82_22# a_82_22# VSUBS a_82_22# m1_126_952#
+ m1_30_110# m1_30_110# a_82_22# a_82_22# m1_30_728# a_82_22# m1_126_952# m1_30_728#
+ m1_30_728# a_82_22# m1_30_110# m1_30_728# a_82_22# a_82_22# m1_30_110# m1_30_728#
+ a_82_22# a_82_22# m1_126_952# a_82_22# a_82_22# a_82_22# a_82_22# a_82_22# m1_30_110#
+ a_82_22# m1_126_952# m1_30_728# m1_30_110# m1_30_728# a_82_22# m1_30_728# m1_30_110#
+ m1_30_728# m1_126_952# a_82_22# m1_30_728# m1_30_110# m1_126_952# a_82_22# a_82_22#
+ a_82_22# a_82_22# a_82_22# a_82_22# a_82_22# m1_30_728# a_82_22# sky130_fd_pr__nfet_01v8_lvt_RE4MKQ
.ends

.subckt sky130_fd_sc_hs__inv_4 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=6.72e+11p pd=5.68e+06u as=9.968e+11p ps=8.5e+06u w=1.12e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=4.44e+11p pd=4.16e+06u as=6.882e+11p ps=6.3e+06u w=740000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG#3 m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ZHX6G9 a_n383_109# a_n29_n509# a_380_21# a_n92_21#
+ a_n682_n597# a_n619_109# a_561_109# a_89_n509# a_n210_n597# a_n564_n597# a_207_109#
+ a_n29_109# a_n501_n509# a_n737_109# a_380_n597# a_n92_n597# a_n446_n597# a_26_21#
+ a_561_n509# a_n147_109# a_n383_n509# a_679_109# a_n328_21# a_n446_21# a_n737_n509#
+ a_n564_21# a_262_n597# a_n328_n597# a_n682_21# a_325_109# a_443_n509# a_616_n597#
+ a_n265_n509# a_n210_21# a_89_109# a_n619_n509# a_144_n597# a_n265_109# a_n839_n683#
+ a_498_n597# a_n501_109# a_325_n509# a_679_n509# a_n147_n509# a_616_21# a_498_21#
+ a_443_109# a_144_21# a_207_n509# a_26_n597# a_262_21#
X0 a_89_109# a_26_21# a_n29_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X1 a_n383_n509# a_n446_n597# a_n501_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X2 a_n147_109# a_n210_21# a_n265_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X3 a_679_109# a_616_21# a_561_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X4 a_n619_n509# a_n682_n597# a_n737_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X5 a_n29_n509# a_n92_n597# a_n147_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X6 a_443_109# a_380_21# a_325_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X7 a_561_109# a_498_21# a_443_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X8 a_325_n509# a_262_n597# a_207_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X9 a_325_109# a_262_21# a_207_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X10 a_n265_n509# a_n328_n597# a_n383_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X11 a_561_n509# a_498_n597# a_443_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X12 a_n619_109# a_n682_21# a_n737_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X13 a_207_109# a_144_21# a_89_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X14 a_n501_109# a_n564_21# a_n619_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X15 a_89_n509# a_26_n597# a_n29_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X16 a_207_n509# a_144_n597# a_89_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 a_n501_n509# a_n564_n597# a_n619_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 a_n147_n509# a_n210_n597# a_n265_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 a_n383_109# a_n446_21# a_n501_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X20 a_679_n509# a_616_n597# a_561_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X21 a_n29_109# a_n92_21# a_n147_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X22 a_n265_109# a_n328_21# a_n383_109# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X23 a_443_n509# a_380_n597# a_325_n509# a_n839_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
.ends

.subckt lvds_diffamp m1_70_160# m1_188_1002# m1_70_80# m1_70_700# m1_188_384# m1_70_778#
+ VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_ZHX6G9_0 m1_188_1002# m1_70_160# m1_70_700# m1_70_700#
+ m1_70_80# m1_188_1002# m1_188_1002# m1_188_384# m1_70_80# m1_70_80# m1_70_778# m1_70_778#
+ m1_70_160# m1_70_778# m1_70_80# m1_70_80# m1_70_80# m1_70_700# m1_188_384# m1_188_1002#
+ m1_188_384# m1_70_778# m1_70_700# m1_70_700# m1_70_160# m1_70_700# m1_70_80# m1_70_80#
+ m1_70_700# m1_188_1002# m1_70_160# m1_70_80# m1_70_160# m1_70_700# m1_188_1002#
+ m1_188_384# m1_70_80# m1_70_778# VSUBS m1_70_80# m1_70_778# m1_188_384# m1_70_160#
+ m1_188_384# m1_70_700# m1_70_700# m1_70_778# m1_70_700# m1_70_160# m1_70_80# m1_70_700#
+ sky130_fd_pr__nfet_01v8_lvt_ZHX6G9
.ends

.subckt transmitter VN m1_20_640# In
Xlvds_currm_n_7 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_26 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_15 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_8 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_27 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_16 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_9 m2_17470_3120# m2_18900_460# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_28 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_17 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_29 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_18 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_19 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xsky130_fd_pr__res_xhigh_po_0p35_ZPVFQL_0 OutN VN m1_13800_6190# vm20g m1_13800_6190#
+ sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL
Xsky130_fd_pr__res_xhigh_po_0p35_ZPVFQL_1 vm20g VN m1_14510_6190# OutP m1_14510_6190#
+ sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL
Xsky130_fd_pr__res_xhigh_po_0p35_ZPVFQL_2 m1_15390_3750# VN VP m1_15390_3750# m1_15690_6180#
+ sky130_fd_pr__res_xhigh_po_0p35_ZPVFQL
Xsky130_fd_sc_hs__inv_16_0 vx9y VN VP vx6y VN VP sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_1 vx6y VN VP vm5g VN VP sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_2 vx6y VN VP vm5g VN VP sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_3 vx6y VN VP vm5g VN VP sky130_fd_sc_hs__inv_16
Xsky130_fd_pr__res_xhigh_po_0p35_RS2YEK_0 m1_16410_6170# m1_16110_3750# m1_16110_3750#
+ m1_16410_6170# VN m1_15690_6180# VN sky130_fd_pr__res_xhigh_po_0p35_RS2YEK
Xsky130_fd_sc_hs__inv_16_4 vx6y VN VP vm5g VN VP sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_5 vx1y VN VP vm2g VN VP sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_6 vx1y VN VP vm2g VN VP sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_7 vx1y VN VP vm2g VN VP sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_8 vx14y VN VP vx1y VN VP sky130_fd_sc_hs__inv_16
Xlvds_currm_p_30 m2_19260_4160# m2_19260_4160# lvds_currm_p_30/m1_60_1070# VP lvds_currm_p
Xsky130_fd_sc_hs__inv_16_9 vx1y VN VP vm2g VN VP sky130_fd_sc_hs__inv_16
Xlvds_currm_p_20 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_22 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_21 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_11 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_10 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_23 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_12 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_switch_p_0 OutN vm6d OutN vm6d OutN vm2g vm6d VP lvds_switch_p
Xlvds_currm_p_24 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_13 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_switch_p_1 OutP vm6d OutP vm6d OutP vm5g vm6d VP lvds_switch_p
Xlvds_currm_p_25 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_14 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_26 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_15 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_27 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_16 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_0 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xsky130_fd_pr__cap_mim_m3_1_N3PKNJ_0 vm20g m1_17940_7520# sky130_fd_pr__cap_mim_m3_1_N3PKNJ
Xlvds_nswitch_0 vm1d OutN OutN vm2g VN lvds_nswitch
Xlvds_currm_p_28 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_17 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_1 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_nswitch_1 vm1d OutP OutP vm5g VN lvds_nswitch
Xlvds_currm_p_29 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_18 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_2 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xsky130_fd_sc_hs__inv_4_0 In VN VP vx9y VN VP sky130_fd_sc_hs__inv_4
Xlvds_currm_p_19 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_3 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_n_0 m1_20_640# lvds_currm_n_0/m1_n20_420# m1_20_640# VN lvds_currm_n
Xsky130_fd_sc_hs__inv_4_1 vx9y VN VP vx14y VN VP sky130_fd_sc_hs__inv_4
Xlvds_currm_n_30 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_p_4 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_0 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#3
Xlvds_currm_n_1 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_31 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_20 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_p_5 m1_17940_7520# m1_17940_7520# m2_17720_10420# VP lvds_currm_p
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_1 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#3
Xlvds_currm_n_10 m2_17470_3120# m2_18900_460# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_2 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_21 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_p_7 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_p_6 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_diffamp_1 m2_17470_3120# m2_17470_3120# m1_15690_6180# m1_15690_6180# m2_19260_4160#
+ m2_19260_4160# VN lvds_diffamp
Xlvds_diffamp_0 m2_17470_3120# m2_17470_3120# vm20g vm20g m1_17940_7520# m1_17940_7520#
+ VN lvds_diffamp
Xlvds_currm_n_11 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_3 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_22 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_p_8 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_n_5 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_4 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_23 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_12 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_p_9 m2_19260_4160# vm6d m3_9390_18600# VP lvds_currm_p
Xlvds_currm_n_6 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_25 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_24 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_14 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
Xlvds_currm_n_13 vm1d m2_1870_1020# m1_20_640# VN lvds_currm_n
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2 m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WXTTNJ c1_n2050_n2000# m3_n2150_n2100#
X0 c1_n2050_n2000# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
.ends

.subckt sky130_fd_pr__res_high_po_5p73_PA2QZX a_n573_400# a_n573_n832# a_n703_n962#
X0 a_n573_n832# a_n573_400# a_n703_n962# sky130_fd_pr__res_high_po_5p73 l=4e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_324MKY a_n369_n509# a_n81_109# a_n129_531# a_303_n509#
+ a_351_n87# a_n33_n87# a_399_109# a_n129_n597# a_n513_n597# a_63_n597# a_n273_109#
+ a_n465_n509# a_n225_n87# a_447_531# a_15_109# a_n321_531# a_15_n509# a_n177_n509#
+ a_111_n509# a_n321_n597# a_207_109# a_n417_n87# a_n465_109# a_n273_n509# a_351_21#
+ a_n513_531# a_n33_21# a_n225_21# a_n177_109# a_447_n597# a_n557_n509# a_495_109#
+ a_399_n509# a_n81_n509# a_111_109# a_n557_109# a_n369_109# a_159_21# a_495_n509#
+ a_63_531# a_255_n597# a_n659_n683# a_159_n87# a_n417_21# a_303_109# a_255_531# a_207_n509#
X0 a_399_n509# a_351_n87# a_303_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n81_109# a_n129_531# a_n177_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_111_109# a_63_531# a_15_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n465_n509# a_n513_n597# a_n557_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X4 a_n273_109# a_n321_531# a_n369_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_n177_109# a_n225_21# a_n273_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 a_n81_n509# a_n129_n597# a_n177_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_15_n509# a_n33_n87# a_n81_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X8 a_n369_n509# a_n417_n87# a_n465_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X9 a_303_n509# a_255_n597# a_207_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_n273_n509# a_n321_n597# a_n369_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_303_109# a_255_531# a_207_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_207_109# a_159_21# a_111_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 a_399_109# a_351_21# a_303_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X14 a_495_109# a_447_531# a_399_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X15 a_n177_n509# a_n225_n87# a_n273_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 a_207_n509# a_159_n87# a_111_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17 a_495_n509# a_447_n597# a_399_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X18 a_n465_109# a_n513_531# a_n557_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X19 a_n369_109# a_n417_21# a_n465_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 a_111_n509# a_63_n597# a_15_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 a_15_109# a_n33_21# a_n81_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt outd_diffamp m1_610_8380# m1_226_8380# m1_802_8758# m1_418_8758# m1_2276_8758#
+ m1_2084_8380# m1_1700_8758# m1_1186_8380# m1_898_8998# m1_130_8998# m1_706_8140#
+ m1_1796_8998# m1_1090_8998# m1_2564_8140# m1_1604_8140# m1_610_8758# m1_226_8758#
+ m1_2084_8758# m1_1186_8758# m1_514_8140# m1_706_8998# m1_2564_8998# m1_2372_8140#
+ m1_1604_8998# m1_994_8380# a_1560_8562# m1_2468_8380# m1_1892_8380# a_182_8562#
+ m1_1508_8380# m1_514_8998# a_1560_9180# m1_322_8140# m1_2180_8140# m1_2372_8998#
+ m1_1988_8140# m1_994_8758# a_182_9180# m1_802_8380# m1_418_8380# m1_1892_8758# VSUBS
+ m1_2276_8380# m1_2468_8758# m1_1700_8380# m1_1508_8758# m1_322_8998# m1_898_8140#
+ m1_130_8140# m1_2180_8998# m1_1796_8140# m1_1090_8140# m1_1988_8998#
Xsky130_fd_pr__nfet_01v8_lvt_324MKY_0 m1_322_8140# m1_610_8758# a_182_9180# m1_994_8380#
+ a_182_8562# a_182_8562# m1_1090_8998# a_182_8562# a_182_8562# a_182_8562# m1_418_8758#
+ m1_226_8380# a_182_8562# a_182_9180# m1_706_8998# a_182_9180# m1_706_8140# m1_514_8140#
+ m1_802_8380# a_182_8562# m1_898_8998# a_182_8562# m1_226_8758# m1_418_8380# a_182_9180#
+ a_182_9180# a_182_9180# a_182_9180# m1_514_8998# a_182_8562# m1_130_8140# m1_1186_8758#
+ m1_1090_8140# m1_610_8380# m1_802_8758# m1_130_8998# m1_322_8998# a_182_9180# m1_1186_8380#
+ a_182_9180# a_182_8562# VSUBS a_182_8562# a_182_9180# m1_994_8758# a_182_9180# m1_898_8140#
+ sky130_fd_pr__nfet_01v8_lvt_324MKY
Xsky130_fd_pr__nfet_01v8_lvt_324MKY_2 m1_2372_8140# m1_2084_8758# a_1560_9180# m1_1700_8380#
+ a_1560_8562# a_1560_8562# m1_1604_8998# a_1560_8562# a_1560_8562# a_1560_8562# m1_2276_8758#
+ m1_2468_8380# a_1560_8562# a_1560_9180# m1_1988_8998# a_1560_9180# m1_1988_8140#
+ m1_2180_8140# m1_1892_8380# a_1560_8562# m1_1796_8998# a_1560_8562# m1_2468_8758#
+ m1_2276_8380# a_1560_9180# a_1560_9180# a_1560_9180# a_1560_9180# m1_2180_8998#
+ a_1560_8562# m1_2564_8140# m1_1508_8758# m1_1604_8140# m1_2084_8380# m1_1892_8758#
+ m1_2564_8998# m1_2372_8998# a_1560_9180# m1_1508_8380# a_1560_9180# a_1560_8562#
+ VSUBS a_1560_8562# a_1560_9180# m1_1700_8758# a_1560_9180# m1_1796_8140# sky130_fd_pr__nfet_01v8_lvt_324MKY
.ends

.subckt sky130_fd_pr__nfet_01v8_ED72KE a_n129_109# a_n753_n1215# a_n753_21# a_n129_727#
+ a_n369_21# a_n705_n509# a_n177_n1215# a_n465_n597# a_255_n509# a_n561_n1215# a_495_n705#
+ a_n609_727# a_n609_109# a_15_1149# a_n273_639# a_399_21# a_n561_1149# a_n81_531#
+ a_447_109# a_447_727# a_399_n1215# a_n177_1149# a_351_n509# a_n417_n509# a_n657_n705#
+ a_n177_n87# a_591_n1215# a_n321_109# a_111_n597# a_n321_727# a_63_n1127# a_n273_531#
+ a_n273_n597# a_n513_n509# a_n797_n1127# a_n33_n1127# a_n129_n509# a_n899_n1301#
+ a_n609_n1127# a_159_109# a_303_n705# a_159_727# a_63_n509# a_n705_n1127# a_n417_n1127#
+ a_n129_n1127# a_n465_639# a_n513_n1127# a_n225_n1127# a_639_727# a_639_109# a_n321_n1127#
+ a_n369_n87# a_n225_n509# a_n465_n705# a_n513_109# a_n513_727# a_687_n597# a_639_n1127#
+ a_n465_531# a_159_n1127# a_447_n1127# a_735_n1127# a_255_n1127# a_543_n1127# a_351_n1127#
+ a_351_727# a_351_109# a_n797_n509# a_n321_n509# a_n33_109# a_n33_727# a_399_1149#
+ a_n81_n597# a_n657_639# a_639_n509# a_111_n705# a_n561_n87# a_n797_727# a_n797_109#
+ a_n225_109# a_n225_727# a_495_639# a_n273_n705# a_15_n1215# a_n705_727# a_n561_21#
+ a_n705_109# a_111_639# a_n177_21# a_n33_n509# a_735_n509# a_n657_531# a_495_n597#
+ a_207_21# a_399_n87# a_543_109# a_543_727# a_591_21# a_495_531# a_111_531# a_591_1149#
+ a_63_727# a_63_109# a_n753_n87# a_n657_n597# a_447_n509# a_687_n705# a_15_n87# a_15_21#
+ a_207_1149# a_n417_109# a_n417_727# a_687_639# a_591_n87# a_303_639# a_n753_1149#
+ a_207_n1215# a_n369_1149# a_255_109# a_255_727# a_543_n509# a_n609_n509# a_159_n509#
+ a_n81_n705# a_207_n87# a_735_727# a_735_109# a_303_n597# a_687_531# a_303_531# a_n369_n1215#
+ a_n81_639#
X0 a_n129_n509# a_n177_n87# a_n225_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n321_n1127# a_n369_n1215# a_n417_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_n417_n509# a_n465_n597# a_n513_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_639_n509# a_591_n87# a_543_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n705_n509# a_n753_n87# a_n797_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X5 a_n33_727# a_n81_639# a_n129_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_351_727# a_303_639# a_255_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_159_727# a_111_639# a_63_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X8 a_255_727# a_207_1149# a_159_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 a_447_727# a_399_1149# a_351_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X10 a_543_727# a_495_639# a_447_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_735_727# a_687_639# a_639_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_63_n1127# a_15_n1215# a_n33_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X13 a_159_n1127# a_111_n705# a_63_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X14 a_639_727# a_591_1149# a_543_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 a_639_n1127# a_591_n1215# a_543_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X16 a_n33_109# a_n81_531# a_n129_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17 a_n33_n509# a_n81_n597# a_n129_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X18 a_351_n509# a_303_n597# a_255_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X19 a_n321_727# a_n369_1149# a_n417_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X20 a_255_n1127# a_207_n1215# a_159_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X21 a_n705_727# a_n753_1149# a_n797_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X22 a_n513_727# a_n561_1149# a_n609_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X23 a_n417_727# a_n465_639# a_n513_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 a_n225_727# a_n273_639# a_n321_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X25 a_n129_727# a_n177_1149# a_n225_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 a_255_109# a_207_21# a_159_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X27 a_351_109# a_303_531# a_255_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X28 a_543_109# a_495_531# a_447_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X29 a_n609_n509# a_n657_n597# a_n705_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X30 a_n417_n1127# a_n465_n705# a_n513_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X31 a_735_n1127# a_687_n705# a_639_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X32 a_n609_727# a_n657_639# a_n705_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 a_159_109# a_111_531# a_63_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X34 a_447_109# a_399_21# a_351_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 a_639_109# a_591_21# a_543_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X36 a_735_109# a_687_531# a_639_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X37 a_n513_n1127# a_n561_n1215# a_n609_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X38 a_351_n1127# a_303_n705# a_255_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X39 a_n513_109# a_n561_21# a_n609_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X40 a_n321_109# a_n369_21# a_n417_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X41 a_n225_109# a_n273_531# a_n321_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X42 a_n705_109# a_n753_21# a_n797_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X43 a_n609_109# a_n657_531# a_n705_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 a_n417_109# a_n465_531# a_n513_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X45 a_n129_109# a_n177_21# a_n225_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 a_255_n509# a_207_n87# a_159_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X47 a_n321_n509# a_n369_n87# a_n417_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X48 a_63_727# a_15_1149# a_n33_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 a_543_n509# a_495_n597# a_447_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X50 a_n33_n1127# a_n81_n705# a_n129_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X51 a_63_109# a_15_21# a_n33_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 a_159_n509# a_111_n597# a_63_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X53 a_n225_n509# a_n273_n597# a_n321_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 a_447_n509# a_399_n87# a_351_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 a_n129_n1127# a_n177_n1215# a_n225_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X56 a_447_n1127# a_399_n1215# a_351_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X57 a_n609_n1127# a_n657_n705# a_n705_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X58 a_n513_n509# a_n561_n87# a_n609_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X59 a_63_n509# a_15_n87# a_n33_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 a_735_n509# a_687_n597# a_639_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X61 a_n225_n1127# a_n273_n705# a_n321_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 a_543_n1127# a_495_n705# a_447_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 a_n705_n1127# a_n753_n1215# a_n797_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_A574RZ a_761_1345# a_1235_109# a_1235_727# a_n1135_727#
+ a_n1135_109# a_n1135_n1127# a_n1135_n1745# a_n977_n2363# a_n29_n509# a_n503_n1127#
+ a_n503_n1745# a_n129_n2451# a_n29_1963# a_29_n597# a_n29_1345# a_977_21# a_n1235_n2451#
+ a_n129_n597# a_187_21# a_n603_n2451# a_n187_n509# a_n345_n1745# a_n603_639# a_n345_n1127#
+ a_187_n597# a_1077_109# a_n977_109# a_1077_727# a_n977_727# a_1135_639# a_n819_n1745#
+ a_n187_1963# a_n819_n1127# a_n187_1345# a_29_n1215# a_29_n1833# a_n1077_n2451# a_503_n2451#
+ a_n445_n2451# a_129_109# a_129_727# a_n187_n1745# a_n445_21# a_29_1257# a_29_1875#
+ a_n187_n1127# a_n919_n2451# a_1135_n2451# a_n1293_n1745# a_n287_n597# a_n129_1875#
+ a_n1293_n1127# a_n819_n509# a_n129_1257# a_n445_639# a_n661_n1745# a_345_n2451#
+ a_819_n597# a_n819_1963# a_n661_n1127# a_n287_n2451# a_977_639# a_n819_1345# a_187_1257#
+ a_187_1875# a_819_n2451# a_n345_n509# a_n1077_n597# a_345_n597# a_n1077_21# a_n345_1345#
+ a_n345_1963# a_n29_727# a_n761_n2451# a_n29_109# a_187_n2451# a_n1135_n509# a_n919_n597#
+ a_345_21# a_29_21# a_n977_n1127# a_n977_n1745# a_n287_1875# a_n977_n509# a_n287_1257#
+ a_n287_639# a_n1135_1345# a_n1135_1963# a_977_n597# a_n503_727# a_n129_n1215# a_n129_n1833#
+ a_129_n2363# a_n445_n597# a_n503_109# a_819_1257# a_n977_1963# a_819_1875# a_661_n2451#
+ a_603_109# a_603_727# a_n977_1345# a_n1235_n1833# a_n1077_1257# a_n1077_1875# a_n1235_n1215#
+ a_29_639# a_345_1875# a_345_1257# a_n603_n1215# a_n603_n1833# a_603_n2363# a_n1235_n597#
+ a_n603_21# a_n503_n509# a_129_n509# a_n1293_n509# a_n1293_109# a_n1293_727# a_1235_n2363#
+ a_503_n597# a_n919_1875# a_977_n2451# a_n503_1345# a_n919_1257# a_n503_1963# a_n1077_n1833#
+ a_n1077_n1215# a_129_1345# a_129_1963# a_n1293_1963# a_n1293_1345# a_n345_727# a_n919_639#
+ a_503_n1215# a_n445_n1833# a_503_n1833# a_445_n2363# a_n345_109# a_977_1257# a_977_1875#
+ a_n445_n1215# a_445_109# a_445_727# a_503_639# a_n445_1257# a_n445_1875# a_n919_n1833#
+ a_919_n2363# a_n919_n1215# a_n1235_21# a_1135_n1215# a_1135_n1833# a_1077_n2363#
+ a_n603_n597# a_1135_n597# a_n661_n509# a_n761_639# a_287_n509# a_n1235_1257# a_n1235_1875#
+ a_345_n1215# a_n287_n1833# a_345_n1833# a_287_n2363# a_661_n597# a_503_21# a_n287_n1215#
+ a_819_n1833# a_n661_1963# a_503_1875# a_819_n1215# a_n661_1345# a_503_1257# a_287_1963#
+ a_287_1345# a_n187_109# a_n187_727# a_287_727# a_n761_n1833# a_761_n2363# a_287_109#
+ a_345_639# a_n761_n1215# a_187_n1833# a_n29_n2363# a_187_n1215# a_n761_n597# a_n603_1257#
+ a_1135_1875# a_n603_1875# a_919_n509# a_1135_1257# a_129_n1745# a_1135_21# a_n1395_n2537#
+ a_129_n1127# a_661_n1833# a_661_n1215# a_n919_21# a_661_1257# a_919_1963# a_661_1875#
+ a_919_1345# a_n761_21# a_445_n509# a_n129_21# a_n819_727# a_603_n1745# a_n819_109#
+ a_187_639# a_603_n1127# a_n1135_n2363# a_919_109# a_919_727# a_445_1963# a_445_1345#
+ a_1235_n1745# a_977_n1215# a_1235_n1127# a_977_n1833# a_n503_n2363# a_n761_1875#
+ a_n761_1257# a_n1235_639# a_n661_109# a_n661_727# a_445_n1745# a_1077_n509# a_761_727#
+ a_445_n1127# a_761_109# a_919_n1127# a_919_n1745# a_819_21# a_1077_1963# a_1077_n1127#
+ a_1077_n1745# a_661_21# a_1077_1345# a_n345_n2363# a_n819_n2363# a_819_639# a_29_n2451#
+ a_287_n1127# a_287_n1745# a_603_n509# a_603_1345# a_603_1963# a_n187_n2363# a_n1077_639#
+ a_661_639# a_761_n1127# a_n29_n1745# a_761_n1745# a_n29_n1127# a_n1293_n2363# a_n129_639#
+ a_n661_n2363# a_1235_n509# a_761_n509# a_1235_1345# a_1235_1963# a_n287_21# a_761_1963#
X0 a_1235_n1745# a_1135_n1833# a_1077_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_n1135_109# a_n1235_21# a_n1293_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2 a_761_n2363# a_661_n2451# a_603_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3 a_n345_n1127# a_n445_n1215# a_n503_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X4 a_n29_1963# a_n129_1875# a_n187_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X5 a_603_1963# a_503_1875# a_445_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X6 a_1235_n509# a_1135_n597# a_1077_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X7 a_n819_727# a_n919_639# a_n977_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X8 a_n1135_n509# a_n1235_n597# a_n1293_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X9 a_n977_1345# a_n1077_1257# a_n1135_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X10 a_603_n1745# a_503_n1833# a_445_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X11 a_n345_727# a_n445_639# a_n503_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X12 a_1077_1345# a_977_1257# a_919_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X13 a_n661_109# a_n761_21# a_n819_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X14 a_n503_1345# a_n603_1257# a_n661_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X15 a_n819_n1127# a_n919_n1215# a_n977_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X16 a_129_109# a_29_21# a_n29_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X17 a_761_n1745# a_661_n1833# a_603_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X18 a_n977_n1127# a_n1077_n1215# a_n1135_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X19 a_1235_1963# a_1135_1875# a_1077_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X20 a_n503_727# a_n603_639# a_n661_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X21 a_n1135_1963# a_n1235_1875# a_n1293_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X22 a_1235_n1127# a_1135_n1215# a_1077_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X23 a_n187_109# a_n287_21# a_n345_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X24 a_n503_n2363# a_n603_n2451# a_n661_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X25 a_n29_1345# a_n129_1257# a_n187_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X26 a_603_1345# a_503_1257# a_445_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X27 a_287_n2363# a_187_n2451# a_129_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X28 a_n29_727# a_n129_639# a_n187_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X29 a_n819_109# a_n919_21# a_n977_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X30 a_603_n1127# a_503_n1215# a_445_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X31 a_n345_109# a_n445_21# a_n503_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X32 a_n661_n2363# a_n761_n2451# a_n819_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X33 a_n503_n1745# a_n603_n1833# a_n661_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X34 a_761_n1127# a_661_n1215# a_603_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X35 a_n1135_n2363# a_n1235_n2451# a_n1293_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X36 a_n503_109# a_n603_21# a_n661_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X37 a_1077_727# a_977_639# a_919_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X38 a_n1135_1345# a_n1235_1257# a_n1293_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X39 a_1235_1345# a_1135_1257# a_1077_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X40 a_287_n1745# a_187_n1833# a_129_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X41 a_n819_n509# a_n919_n597# a_n977_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X42 a_n661_n1745# a_n761_n1833# a_n819_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X43 a_n29_109# a_n129_21# a_n187_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X44 a_n661_n509# a_n761_n597# a_n819_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X45 a_n29_n2363# a_n129_n2451# a_n187_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X46 a_761_727# a_661_639# a_603_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X47 a_n1135_n1745# a_n1235_n1833# a_n1293_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X48 a_n819_1963# a_n919_1875# a_n977_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X49 a_919_n509# a_819_n597# a_761_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X50 a_n187_n2363# a_n287_n2451# a_n345_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X51 a_n503_n1127# a_n603_n1215# a_n661_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X52 a_287_727# a_187_639# a_129_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X53 a_761_n509# a_661_n597# a_603_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X54 a_1077_109# a_977_21# a_919_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X55 a_n661_1963# a_n761_1875# a_n819_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X56 a_n187_n509# a_n287_n597# a_n345_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X57 a_1235_727# a_1135_639# a_1077_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X58 a_287_n1127# a_187_n1215# a_129_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X59 a_n29_n1745# a_n129_n1833# a_n187_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X60 a_n661_n1127# a_n761_n1215# a_n819_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X61 a_919_727# a_819_639# a_761_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X62 a_919_1963# a_819_1875# a_761_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X63 a_445_727# a_345_639# a_287_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X64 a_n187_n1745# a_n287_n1833# a_n345_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X65 a_n187_1963# a_n287_1875# a_n345_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X66 a_761_1963# a_661_1875# a_603_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X67 a_287_n509# a_187_n597# a_129_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X68 a_761_109# a_661_21# a_603_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X69 a_129_n2363# a_29_n2451# a_n29_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X70 a_n1135_n1127# a_n1235_n1215# a_n1293_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X71 a_n819_1345# a_n919_1257# a_n977_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X72 a_603_727# a_503_639# a_445_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X73 a_287_109# a_187_21# a_129_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X74 a_n661_1345# a_n761_1257# a_n819_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X75 a_1235_109# a_1135_21# a_1077_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X76 a_445_n2363# a_345_n2451# a_287_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X77 a_n29_n1127# a_n129_n1215# a_n187_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X78 a_287_1963# a_187_1875# a_129_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X79 a_129_n1745# a_29_n1833# a_n29_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X80 a_919_1345# a_819_1257# a_761_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X81 a_919_109# a_819_21# a_761_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X82 a_445_109# a_345_21# a_287_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X83 a_n187_n1127# a_n287_n1215# a_n345_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X84 a_n345_n509# a_n445_n597# a_n503_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X85 a_n187_1345# a_n287_1257# a_n345_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X86 a_761_1345# a_661_1257# a_603_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X87 a_919_n2363# a_819_n2451# a_761_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X88 a_445_n1745# a_345_n1833# a_287_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X89 a_129_n509# a_29_n597# a_n29_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X90 a_603_109# a_503_21# a_445_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X91 a_1077_n2363# a_977_n2451# a_919_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X92 a_445_n509# a_345_n597# a_287_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X93 a_n345_1963# a_n445_1875# a_n503_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X94 a_287_1345# a_187_1257# a_129_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X95 a_129_n1127# a_29_n1215# a_n29_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X96 a_919_n1745# a_819_n1833# a_761_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X97 a_129_1963# a_29_1875# a_n29_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X98 a_n345_n2363# a_n445_n2451# a_n503_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X99 a_n977_727# a_n1077_639# a_n1135_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X100 a_1077_n1745# a_977_n1833# a_919_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X101 a_445_1963# a_345_1875# a_287_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X102 a_445_n1127# a_345_n1215# a_287_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X103 a_n977_n509# a_n1077_n597# a_n1135_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X104 a_1077_n509# a_977_n597# a_919_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X105 a_n1135_727# a_n1235_639# a_n1293_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X106 a_n819_n2363# a_n919_n2451# a_n977_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X107 a_n345_1345# a_n445_1257# a_n503_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X108 a_n503_n509# a_n603_n597# a_n661_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X109 a_n345_n1745# a_n445_n1833# a_n503_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X110 a_n977_n2363# a_n1077_n2451# a_n1135_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X111 a_919_n1127# a_819_n1215# a_761_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X112 a_1235_n2363# a_1135_n2451# a_1077_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X113 a_n977_1963# a_n1077_1875# a_n1135_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X114 a_129_1345# a_29_1257# a_n29_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X115 a_n977_109# a_n1077_21# a_n1135_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X116 a_1077_1963# a_977_1875# a_919_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X117 a_n661_727# a_n761_639# a_n819_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X118 a_n503_1963# a_n603_1875# a_n661_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X119 a_1077_n1127# a_977_n1215# a_919_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X120 a_603_n509# a_503_n597# a_445_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X121 a_n29_n509# a_n129_n597# a_n187_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X122 a_445_1345# a_345_1257# a_287_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X123 a_n819_n1745# a_n919_n1833# a_n977_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X124 a_129_727# a_29_639# a_n29_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X125 a_603_n2363# a_503_n2451# a_445_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X126 a_n977_n1745# a_n1077_n1833# a_n1135_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X127 a_n187_727# a_n287_639# a_n345_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
.ends

.subckt outd_cmirror_transistors sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n1745# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n2363#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_1345#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n2363#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_21#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n597#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_1257# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n1745#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_1875#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n2363# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_1345# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n2451#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n2451#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n2451#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_1963#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_1345# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n1833# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_1875#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_1875# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_1875# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n1127#
+ a_2_2306# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n2363#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_1963#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n1215# a_2_1688# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_109# a_2_n58# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_1875#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_1345#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_1257# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n1833#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n597# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n1745# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_639#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n2363#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_n509#
+ VSUBS a_2_560# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n1833#
Xsky130_fd_pr__nfet_01v8_ED72KE_0 sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_109# a_2_n58#
+ a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_727# a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_n509#
+ a_2_n58# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_n509# a_2_n58# a_2_n58#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_109#
+ a_2_2306# a_2_2306# a_2_1688# a_2_2306# a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_727# a_2_n58# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_n509# a_2_n58# a_2_560# a_2_n58# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_109#
+ a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_n1127#
+ a_2_1688# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_n509#
+ VSUBS sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_109#
+ a_2_n58# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_n1127# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_n1127#
+ a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_n509# a_2_n58# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_727# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_n1127#
+ a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_727#
+ a_2_2306# a_2_560# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_n509# a_2_n58#
+ a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_727#
+ a_2_2306# a_2_n58# a_2_n58# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_727# a_2_1688#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_109# a_2_2306# a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_n509# a_2_1688# a_2_560# a_2_1688# a_2_560#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_727#
+ a_2_1688# a_2_1688# a_2_1688# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_109# a_2_560# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_n509#
+ a_2_n58# a_2_560# a_2_1688# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_727# a_2_2306# a_2_560# a_2_2306# a_2_2306#
+ a_2_n58# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_n509# a_2_n58# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_109# a_2_560# a_2_1688# a_2_1688# a_2_n58#
+ a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE
Xsky130_fd_pr__nfet_01v8_A574RZ_0 sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_21# VSUBS sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ
.ends

.subckt outd_cmirror_64t m1_220_5610# m1_0_80# m1_130_5370# VSUBS
Xoutd_cmirror_transistors_0 m1_220_5610# m1_130_5370# m1_130_5370# m1_220_5610# m1_130_5370#
+ VSUBS m1_130_5370# VSUBS m1_220_5610# VSUBS m1_0_80# m1_0_80# VSUBS VSUBS VSUBS
+ m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_220_5610# m1_130_5370# m1_220_5610# m1_220_5610#
+ m1_220_5610# m1_0_80# m1_220_5610# m1_130_5370# m1_220_5610# m1_220_5610# m1_220_5610#
+ VSUBS VSUBS m1_220_5610# VSUBS m1_220_5610# m1_0_80# VSUBS VSUBS m1_0_80# m1_0_80#
+ m1_220_5610# m1_0_80# m1_130_5370# m1_220_5610# m1_220_5610# m1_220_5610# m1_0_80#
+ m1_220_5610# m1_0_80# m1_220_5610# m1_220_5610# m1_220_5610# m1_0_80# m1_220_5610#
+ m1_0_80# m1_220_5610# m1_220_5610# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# VSUBS
+ VSUBS VSUBS m1_130_5370# m1_220_5610# m1_130_5370# VSUBS VSUBS m1_220_5610# m1_0_80#
+ VSUBS VSUBS m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_130_5370# m1_0_80# VSUBS
+ VSUBS m1_220_5610# m1_130_5370# VSUBS m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610#
+ m1_0_80# m1_0_80# VSUBS VSUBS m1_0_80# VSUBS VSUBS m1_220_5610# m1_220_5610# m1_220_5610#
+ m1_130_5370# m1_220_5610# m1_130_5370# m1_130_5370# m1_220_5610# m1_220_5610# m1_0_80#
+ m1_130_5370# m1_220_5610# m1_220_5610# VSUBS VSUBS VSUBS m1_220_5610# m1_220_5610#
+ m1_220_5610# m1_130_5370# m1_220_5610# m1_0_80# m1_130_5370# m1_220_5610# m1_0_80#
+ m1_0_80# VSUBS m1_130_5370# VSUBS VSUBS m1_130_5370# m1_220_5610# m1_220_5610# m1_0_80#
+ m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_220_5610# m1_220_5610# m1_0_80# VSUBS
+ m1_220_5610# m1_0_80# VSUBS m1_0_80# m1_0_80# VSUBS VSUBS m1_220_5610# m1_0_80#
+ m1_0_80# m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS VSUBS m1_0_80# m1_0_80# m1_220_5610#
+ m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS m1_220_5610#
+ VSUBS m1_220_5610# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS
+ m1_220_5610# m1_130_5370# m1_130_5370# m1_0_80# VSUBS VSUBS VSUBS VSUBS m1_220_5610#
+ m1_0_80# m1_220_5610# m1_130_5370# m1_0_80# m1_130_5370# m1_0_80# m1_220_5610# m1_0_80#
+ VSUBS m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_220_5610# m1_220_5610# m1_0_80# m1_0_80#
+ m1_0_80# m1_0_80# m1_0_80# m1_130_5370# m1_130_5370# m1_130_5370# m1_0_80# m1_0_80#
+ m1_0_80# m1_0_80# m1_0_80# m1_130_5370# m1_0_80# m1_0_80# m1_220_5610# m1_220_5610#
+ m1_220_5610# VSUBS m1_220_5610# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_0_80#
+ VSUBS m1_220_5610# m1_0_80# m1_0_80# VSUBS m1_220_5610# VSUBS m1_0_80# m1_0_80#
+ VSUBS VSUBS m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80#
+ m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_220_5610#
+ m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_0_80#
+ m1_220_5610# m1_220_5610# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS m1_220_5610#
+ m1_130_5370# m1_130_5370# m1_220_5610# m1_0_80# m1_0_80# m1_130_5370# m1_130_5370#
+ m1_220_5610# m1_0_80# m1_0_80# m1_130_5370# m1_0_80# m1_0_80# m1_130_5370# VSUBS
+ m1_220_5610# m1_220_5610# VSUBS VSUBS m1_130_5370# m1_0_80# VSUBS m1_0_80# VSUBS
+ m1_0_80# VSUBS m1_130_5370# m1_0_80# m1_130_5370# m1_220_5610# m1_0_80# m1_220_5610#
+ VSUBS VSUBS m1_0_80# VSUBS VSUBS m1_220_5610# m1_0_80# m1_220_5610# m1_0_80# m1_0_80#
+ VSUBS m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS VSUBS VSUBS VSUBS m1_220_5610# m1_220_5610#
+ m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610#
+ VSUBS m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_0_80# outd_cmirror_transistors
.ends

.subckt outd_stage2 m1_370_11400# m1_2350_11400# outd_cmirror_64t_4/m1_0_80# dw_60_8030#
+ m1_1850_8370# m2_7240_7300# cmirror_out m1_250_8900# VN
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_0 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_1 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_2 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_3 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_4 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_5 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_6 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_8 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_7 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_9 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_10 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_11 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_12 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_13 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_14 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_15 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xoutd_diffamp_0 cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_370_11400# m1_2350_11400# m1_2350_11400# cmirror_out cmirror_out cmirror_out
+ cmirror_out m1_370_11400# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400#
+ cmirror_out m1_1850_8370# cmirror_out cmirror_out m1_250_8900# cmirror_out m1_370_11400#
+ m1_1850_8370# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400# cmirror_out
+ m1_250_8900# cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_2350_11400# m1_370_11400# m1_2350_11400# outd_diffamp
Xoutd_cmirror_64t_0 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
Xoutd_diffamp_1 cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_370_11400# m1_2350_11400# m1_2350_11400# cmirror_out cmirror_out cmirror_out
+ cmirror_out m1_370_11400# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400#
+ cmirror_out m1_1850_8370# cmirror_out cmirror_out m1_250_8900# cmirror_out m1_370_11400#
+ m1_1850_8370# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400# cmirror_out
+ m1_250_8900# cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_2350_11400# m1_370_11400# m1_2350_11400# outd_diffamp
Xoutd_cmirror_64t_2 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
Xoutd_cmirror_64t_1 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
Xoutd_diffamp_2 cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_370_11400# m1_2350_11400# m1_2350_11400# cmirror_out cmirror_out cmirror_out
+ cmirror_out m1_370_11400# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400#
+ cmirror_out m1_1850_8370# cmirror_out cmirror_out m1_250_8900# cmirror_out m1_370_11400#
+ m1_1850_8370# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400# cmirror_out
+ m1_250_8900# cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_2350_11400# m1_370_11400# m1_2350_11400# outd_diffamp
Xoutd_cmirror_64t_3 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
Xoutd_diffamp_3 cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_370_11400# m1_2350_11400# m1_2350_11400# cmirror_out cmirror_out cmirror_out
+ cmirror_out m1_370_11400# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400#
+ cmirror_out m1_1850_8370# cmirror_out cmirror_out m1_250_8900# cmirror_out m1_370_11400#
+ m1_1850_8370# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400# cmirror_out
+ m1_250_8900# cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_2350_11400# m1_370_11400# m1_2350_11400# outd_diffamp
Xoutd_cmirror_64t_4 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
.ends

.subckt sky130_fd_pr__nfet_01v8_DJG2KN a_n29_n509# a_29_n597# a_n187_n509# a_n129_n597#
+ a_129_109# a_n289_n683# a_n29_109# a_29_21# a_129_n509# a_n187_109# a_n129_21#
X0 a_129_109# a_29_21# a_n29_109# a_n289_n683# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_n29_109# a_n129_21# a_n187_109# a_n289_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2 a_129_n509# a_29_n597# a_n29_n509# a_n289_n683# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3 a_n29_n509# a_n129_n597# a_n187_n509# a_n289_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt outd_stage3 m4_40470_12200# m3_11690_14240# m2_40400_9110# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ outd_stage2_3/cmirror_out m4_40470_12880# m2_40400_10380# VSUBS
Xoutd_stage2_0 m4_40470_12880# m4_40470_12200# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ m3_11690_14240# m2_40400_9110# m2_41490_8160# outd_stage2_3/cmirror_out m2_40400_10380#
+ VSUBS outd_stage2
Xoutd_stage2_1 m4_40470_12880# m4_40470_12200# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ m3_11690_14240# m2_40400_9110# m2_41490_8160# outd_stage2_3/cmirror_out m2_40400_10380#
+ VSUBS outd_stage2
Xoutd_stage2_2 m4_40470_12880# m4_40470_12200# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ m3_11690_14240# m2_40400_9110# m2_41490_8160# outd_stage2_3/cmirror_out m2_40400_10380#
+ VSUBS outd_stage2
Xoutd_stage2_3 m4_40470_12880# m4_40470_12200# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ m3_11690_14240# m2_40400_9110# m2_41490_8160# outd_stage2_3/cmirror_out m2_40400_10380#
+ VSUBS outd_stage2
.ends

.subckt sky130_fd_pr__nfet_01v8_LH2JGW a_n81_n288# a_63_n200# a_n33_n200# a_15_222#
+ a_n227_n374# a_n125_n200#
X0 a_n33_n200# a_n81_n288# a_n125_n200# a_n227_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X1 a_63_n200# a_15_222# a_n33_n200# a_n227_n374# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__res_high_po_2p85_8GE2XM a_n1512_n1032# a_n694_n1032# a_124_n1032#
+ a_n1512_600# a_n1642_n1162# a_942_n1032# a_124_600# a_942_600# a_n694_600#
X0 a_n1512_n1032# a_n1512_600# a_n1642_n1162# sky130_fd_pr__res_high_po_2p85 l=6e+06u
X1 a_n694_n1032# a_n694_600# a_n1642_n1162# sky130_fd_pr__res_high_po_2p85 l=6e+06u
X2 a_942_n1032# a_942_600# a_n1642_n1162# sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3 a_124_n1032# a_124_600# a_n1642_n1162# sky130_fd_pr__res_high_po_2p85 l=6e+06u
.ends

.subckt outd_stage1 outd_cmirror_64t_0/m1_0_80# m1_n1500_10180# m1_1860_8350# isource_out
+ m1_1830_10170# m1_260_8900# dw_70_8020# VN
Xoutd_cmirror_64t_0 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out
+ VN outd_cmirror_64t
Xoutd_diffamp_0 isource_out isource_out isource_out isource_out isource_out isource_out
+ isource_out isource_out m1_n1500_10180# m1_n1500_10180# m1_n1500_10180# m1_1830_10170#
+ m1_n1500_10180# m1_1830_10170# m1_1830_10170# isource_out isource_out isource_out
+ isource_out m1_n1500_10180# m1_n1500_10180# m1_1830_10170# m1_1830_10170# m1_1830_10170#
+ isource_out m1_1860_8350# isource_out isource_out m1_260_8900# isource_out m1_n1500_10180#
+ m1_1860_8350# m1_n1500_10180# m1_1830_10170# m1_1830_10170# m1_1830_10170# isource_out
+ m1_260_8900# isource_out isource_out isource_out isource_out isource_out isource_out
+ isource_out isource_out m1_n1500_10180# m1_n1500_10180# m1_n1500_10180# m1_1830_10170#
+ m1_1830_10170# m1_n1500_10180# m1_1830_10170# outd_diffamp
Xsky130_fd_pr__res_high_po_2p85_8GE2XM_0 m1_n1500_10180# m1_n1500_10180# m1_n1500_10180#
+ dw_70_8020# VN m1_n1500_10180# dw_70_8020# dw_70_8020# dw_70_8020# sky130_fd_pr__res_high_po_2p85_8GE2XM
Xsky130_fd_pr__res_high_po_2p85_8GE2XM_1 m1_1830_10170# m1_1830_10170# m1_1830_10170#
+ dw_70_8020# VN m1_1830_10170# dw_70_8020# dw_70_8020# dw_70_8020# sky130_fd_pr__res_high_po_2p85_8GE2XM
.ends

.subckt outd VP InputRef I_Bias outd_stage1_0/isource_out VM1_D VM14D InputSignal
+ VN
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_6 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_7 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_1_WXTTNJ_0 VN I_Bias sky130_fd_pr__cap_mim_m3_1_WXTTNJ
Xsky130_fd_pr__cap_mim_m3_1_WXTTNJ_1 VN I_Bias sky130_fd_pr__cap_mim_m3_1_WXTTNJ
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_8 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xoutd_stage2_0 V_da2_N V_da2_P I_Bias VP V_da1_P outd_stage2_0/m2_7240_7300# VM1_D
+ V_da1_N VN outd_stage2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_9 VN InputRef sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__nfet_01v8_DJG2KN_0 m1_n19890_7120# I_Bias VN I_Bias VN VN m1_n19890_7120#
+ I_Bias VN VN I_Bias sky130_fd_pr__nfet_01v8_DJG2KN
Xoutd_stage3_0 OutputP VP V_da2_P I_Bias VM14D OutputN V_da2_N VN outd_stage3
Xsky130_fd_pr__nfet_01v8_LH2JGW_0 I_Bias m1_n19890_7120# I_Bias I_Bias VN m1_n19890_7120#
+ sky130_fd_pr__nfet_01v8_LH2JGW
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_10 VN InputRef sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xoutd_stage1_0 I_Bias V_da1_P InputRef outd_stage1_0/isource_out V_da1_N InputSignal
+ VP VN outd_stage1
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_0 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_1 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_2 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_4 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_3 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_5 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
.ends

.subckt sky130_fd_pr__nfet_01v8_6YE2KS a_n345_n200# a_129_n200# a_287_n200# a_29_n288#
+ a_n129_n288# a_187_n288# a_n287_n288# a_n29_n200# a_n187_n200# a_n447_n374#
X0 a_n187_n200# a_n287_n288# a_n345_n200# a_n447_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_287_n200# a_187_n288# a_129_n200# a_n447_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2 a_129_n200# a_29_n288# a_n29_n200# a_n447_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3 a_n29_n200# a_n129_n288# a_n187_n200# a_n447_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_QQ8PGA a_255_n509# a_n129_109# a_15_n597# a_111_21#
+ a_351_n509# a_n177_n597# a_n321_109# a_n515_n683# a_n129_n509# a_111_n87# a_15_531#
+ a_63_n509# a_159_109# a_n225_n509# a_207_531# a_n81_21# a_n273_21# a_n321_n509#
+ a_351_109# a_n33_109# a_303_21# a_303_n87# a_n225_109# a_n413_109# a_n177_531# a_n33_n509#
+ a_n81_n87# a_n273_n87# a_63_109# a_207_n597# a_n369_531# a_159_n509# a_n369_n597#
+ a_255_109# a_n413_n509#
X0 a_n129_n509# a_n177_n597# a_n225_n509# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n33_109# a_n81_21# a_n129_109# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_n33_n509# a_n81_n87# a_n129_n509# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X3 a_351_n509# a_303_n87# a_255_n509# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_255_109# a_207_531# a_159_109# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_351_109# a_303_21# a_255_109# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X6 a_159_109# a_111_21# a_63_109# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_n321_109# a_n369_531# a_n413_109# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X8 a_n225_109# a_n273_21# a_n321_109# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X9 a_n129_109# a_n177_531# a_n225_109# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 a_255_n509# a_207_n597# a_159_n509# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X11 a_n321_n509# a_n369_n597# a_n413_n509# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X12 a_63_109# a_15_531# a_n33_109# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 a_159_n509# a_111_n87# a_63_n509# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X14 a_n225_n509# a_n273_n87# a_n321_n509# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 a_63_n509# a_15_n597# a_n33_n509# a_n515_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt bias_curm_n m1_80_970# m1_176_1194# a_132_882# VSUBS
Xsky130_fd_pr__nfet_01v8_6YE2KS_0 VSUBS m1_80_970# VSUBS a_132_882# a_132_882# a_132_882#
+ a_132_882# VSUBS m1_80_970# VSUBS sky130_fd_pr__nfet_01v8_6YE2KS
Xsky130_fd_pr__nfet_01v8_QQ8PGA_0 m1_176_1194# m1_176_1194# a_132_882# a_132_882#
+ m1_80_970# a_132_882# m1_176_1194# VSUBS m1_176_1194# a_132_882# a_132_882# m1_176_1194#
+ m1_80_970# m1_80_970# a_132_882# a_132_882# a_132_882# m1_176_1194# m1_80_970# m1_80_970#
+ a_132_882# a_132_882# m1_80_970# m1_80_970# a_132_882# m1_80_970# a_132_882# a_132_882#
+ m1_176_1194# a_132_882# a_132_882# m1_80_970# a_132_882# m1_176_1194# m1_80_970#
+ sky130_fd_pr__nfet_01v8_QQ8PGA
.ends

.subckt eight-mirrors-p m3_590_440# m2_150_1940# m1_910_120#
Xbias_curm_p_6 m3_590_440# m2_920_6270# m1_910_120# m2_150_1940# bias_curm_p
Xbias_curm_p_7 m3_590_440# m2_920_6270# m1_910_120# m2_150_1940# bias_curm_p
Xbias_curm_p_0 m3_590_440# m2_920_6270# m1_910_120# m2_150_1940# bias_curm_p
Xbias_curm_p_1 m3_590_440# m2_920_6270# m1_910_120# m2_150_1940# bias_curm_p
Xbias_curm_p_2 m3_590_440# m2_920_6270# m1_910_120# m2_150_1940# bias_curm_p
Xbias_curm_p_3 m3_590_440# m2_920_6270# m1_910_120# m2_150_1940# bias_curm_p
Xbias_curm_p_4 m3_590_440# m2_920_6270# m1_910_120# m2_150_1940# bias_curm_p
Xbias_curm_p_5 m3_590_440# m2_920_6270# m1_910_120# m2_150_1940# bias_curm_p
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_26U9NK c2_n3251_n1500# m4_n3351_n1600#
X0 c2_n3251_n1500# m4_n3351_n1600# sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt curr_mirror_channel TIA_Bias Comp_Bias_6 Comp_Bias_5 ctl_Bias VP Comp_Bias_3
+ Comp_Bias_2 Comp_Bias_1 LVDS_Bias I_in m3_14070_2720# Bias_Analog_out VSUBS
Xbias_curm_p_6 TIA_Bias m2_3110_8460# vm12d VP bias_curm_p
Xbias_curm_n_3 m2_3220_480# vm12d I_in VSUBS bias_curm_n
Xbias_curm_p_7 FB_Bias_1 bias_curm_p_7/m1_120_n692# vm4d VP bias_curm_p
Xbias_curm_p_8 ctl_Bias m2_6380_8570# vm12d VP bias_curm_p
Xbias_curm_p_9 Bias_Analog_out m2_5290_6250# vm12d VP bias_curm_p
Xbias_curm_p_10 Bias_Analog_out m2_5290_6250# vm12d VP bias_curm_p
Xbias_curm_p_11 Bias_Analog_out m2_5290_6250# vm12d VP bias_curm_p
Xbias_curm_p_12 ctl_Bias m2_6380_8570# vm12d VP bias_curm_p
Xbias_curm_p_13 Bias_Analog_out m2_5290_6250# vm12d VP bias_curm_p
Xbias_curm_p_14 Bias_Analog_out m2_5290_6250# vm12d VP bias_curm_p
Xbias_curm_p_15 Bias_Analog_out m2_5290_6250# vm12d VP bias_curm_p
Xbias_curm_p_16 ctl_Bias m2_6380_8570# vm12d VP bias_curm_p
Xbias_curm_p_17 ctl_Bias m2_6380_8570# vm12d VP bias_curm_p
Xeight-mirrors-p_0 Comp_Bias_1 VP vm12d eight-mirrors-p
Xeight-mirrors-p_1 Comp_Bias_2 VP vm12d eight-mirrors-p
Xeight-mirrors-p_2 m3_14070_2720# VP vm12d eight-mirrors-p
Xeight-mirrors-p_3 Comp_Bias_3 VP vm12d eight-mirrors-p
Xeight-mirrors-p_4 Comp_Bias_6 VP vm12d eight-mirrors-p
Xsky130_fd_pr__cap_mim_m3_2_26U9NK_0 VP vm4d sky130_fd_pr__cap_mim_m3_2_26U9NK
Xeight-mirrors-p_5 Comp_Bias_5 VP vm12d eight-mirrors-p
Xsky130_fd_pr__cap_mim_m3_2_26U9NK_1 VP vm12d sky130_fd_pr__cap_mim_m3_2_26U9NK
Xeight-mirrors-p_6 LVDS_Bias VP vm12d eight-mirrors-p
Xbias_curm_p_0 vm4d bias_curm_p_0/m1_120_n692# vm4d VP bias_curm_p
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_1 VSUBS VP sky130_fd_pr__cap_mim_m3_2_LJ5JLG
Xbias_curm_p_1 vm12d bias_curm_p_1/m1_120_n692# vm12d VP bias_curm_p
Xbias_curm_p_3 TIA_Bias m2_3110_8460# vm12d VP bias_curm_p
Xbias_curm_p_2 TIA_Bias m2_3110_8460# vm12d VP bias_curm_p
Xbias_curm_p_4 TIA_Bias m2_3110_8460# vm12d VP bias_curm_p
Xbias_curm_n_1 bias_curm_n_1/m1_80_970# vm4d I_in VSUBS bias_curm_n
Xbias_curm_n_0 bias_curm_n_0/m1_80_970# I_in I_in VSUBS bias_curm_n
Xbias_curm_p_5 TIA_Bias m2_3110_8460# vm12d VP bias_curm_p
Xbias_curm_n_2 m2_3220_480# vm12d I_in VSUBS bias_curm_n
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL a_n642_n1562# a_442_1000# a_n194_n1432#
+ a_n194_1000# a_442_n1432# a_n512_n1432# a_124_n1432# a_n512_1000# a_124_1000#
X0 a_n512_n1432# a_n512_1000# a_n642_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
X1 a_124_n1432# a_124_1000# a_n642_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
X2 a_n194_n1432# a_n194_1000# a_n642_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
X3 a_442_n1432# a_442_1000# a_n642_n1562# sky130_fd_pr__res_xhigh_po_0p35 l=1e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_HR8DH9 a_262_n288# a_n328_n288# a_n501_n200# a_616_n288#
+ a_561_n200# a_144_n288# a_n839_n374# a_n383_n200# a_498_n288# a_n737_n200# a_443_n200#
+ a_n265_n200# a_n619_n200# a_26_n288# a_325_n200# a_n682_n288# a_679_n200# a_n147_n200#
+ a_207_n200# a_n210_n288# a_n564_n288# a_n29_n200# a_380_n288# a_n92_n288# a_89_n200#
+ a_n446_n288#
X0 a_325_n200# a_262_n288# a_207_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X1 a_n265_n200# a_n328_n288# a_n383_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X2 a_561_n200# a_498_n288# a_443_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X3 a_89_n200# a_26_n288# a_n29_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X4 a_207_n200# a_144_n288# a_89_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X5 a_n501_n200# a_n564_n288# a_n619_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X6 a_n147_n200# a_n210_n288# a_n265_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X7 a_679_n200# a_616_n288# a_561_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X8 a_443_n200# a_380_n288# a_325_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X9 a_n383_n200# a_n446_n288# a_n501_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10 a_n619_n200# a_n682_n288# a_n737_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X11 a_n29_n200# a_n92_n288# a_n147_n200# a_n839_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
.ends

.subckt currm_comp m1_522_170# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n328_n288# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_498_n288#
+ m1_994_170# m1_50_170# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_26_n288# m1_1230_170#
+ m1_1348_410# m1_168_410# m1_404_410# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n682_n288#
+ m1_758_170# m1_876_410# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n210_n288# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n92_n288#
+ sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_380_n288# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n564_n288#
+ m1_1112_410# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n446_n288# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_262_n288#
+ m1_1466_170# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_616_n288# m1_286_170# m1_640_410#
+ VSUBS sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_144_n288#
Xsky130_fd_pr__nfet_01v8_lvt_HR8DH9_0 sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_262_n288#
+ sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n328_n288# m1_286_170# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_616_n288#
+ m1_1348_410# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_144_n288# VSUBS m1_404_410#
+ sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_498_n288# m1_50_170# m1_1230_170# m1_522_170#
+ m1_168_410# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_26_n288# m1_1112_410# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n682_n288#
+ m1_1466_170# m1_640_410# m1_994_170# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n210_n288#
+ sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n564_n288# m1_758_170# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_380_n288#
+ sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n92_n288# m1_876_410# sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0/a_n446_n288#
+ sky130_fd_pr__nfet_01v8_lvt_HR8DH9
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_DG2JGC a_15_n200# a_n177_n200# a_111_n200# a_n273_n200#
+ a_159_n288# a_63_222# a_n81_n200# a_255_222# a_399_n200# a_351_n288# a_n417_n288#
+ a_n129_222# a_n563_n374# a_207_n200# a_n225_n288# a_n321_222# a_n461_n200# a_n369_n200#
+ a_303_n200# a_n33_n288#
X0 a_n81_n200# a_n129_222# a_n177_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_15_n200# a_n33_n288# a_n81_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X2 a_n369_n200# a_n417_n288# a_n461_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X3 a_303_n200# a_255_222# a_207_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n273_n200# a_n321_222# a_n369_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X5 a_207_n200# a_159_n288# a_111_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_n177_n200# a_n225_n288# a_n273_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 a_111_n200# a_63_222# a_15_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 a_399_n200# a_351_n288# a_303_n200# a_n563_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt diffamp_element m1_838_660# m1_934_420# a_698_850# m1_646_660# a_890_840#
+ VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_DG2JGC_0 m1_838_660# m1_838_660# m1_934_420# VSUBS a_890_840#
+ a_890_840# m1_934_420# a_890_840# m1_838_660# a_890_840# VSUBS a_890_840# VSUBS
+ m1_838_660# a_698_850# a_698_850# VSUBS m1_646_660# m1_934_420# a_890_840# sky130_fd_pr__nfet_01v8_lvt_DG2JGC
.ends

.subckt sky130_fd_pr__res_xhigh_po_2p85_TY94YJ a_n285_100# a_n285_n532# a_n415_n662#
X0 a_n285_n532# a_n285_100# a_n415_n662# sky130_fd_pr__res_xhigh_po_2p85 l=1e+06u
.ends

.subckt comp_adv3_di Outn bias VP diffamp_element_0/a_890_840# diffamp_element_1/a_890_840#
+ Outp VN
Xcurrm_comp_0 VN bias bias VN VN bias VN m2_820_n490# bias m2_820_n490# VN VN m2_820_n490#
+ bias bias bias bias m2_820_n490# bias bias VN bias VN m2_820_n490# VN bias currm_comp
Xdiffamp_element_0 Outp m2_820_n490# Inn2 Inn2 diffamp_element_0/a_890_840# VN diffamp_element
Xdiffamp_element_1 Outn m2_820_n490# Inp2 Inp2 diffamp_element_1/a_890_840# VN diffamp_element
Xsky130_fd_pr__res_xhigh_po_2p85_TY94YJ_0 VP Outn VN sky130_fd_pr__res_xhigh_po_2p85_TY94YJ
Xsky130_fd_pr__res_xhigh_po_2p85_TY94YJ_1 VP Outp VN sky130_fd_pr__res_xhigh_po_2p85_TY94YJ
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_MJMGTW c2_n3251_n2000# m4_n3351_n2100#
X0 c2_n3251_n2000# m4_n3351_n2100# sky130_fd_pr__cap_mim_m3_2 l=2e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_H9XL9H c1_n550_n500# m3_n650_n600#
X0 c1_n550_n500# m3_n650_n600# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_2p85_8K9944 a_n285_150# a_n285_n582# a_n415_n712#
X0 a_n285_n582# a_n285_150# a_n415_n712# sky130_fd_pr__res_xhigh_po_2p85 l=1.5e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_V6SMGN a_n129_n200# a_n81_n288# a_63_n200# a_n177_222#
+ a_n225_n200# a_n33_n200# a_n419_n374# a_n317_n200# a_159_n200# a_111_n288# a_15_222#
+ a_n273_n288# a_255_n200# a_207_222#
X0 a_n33_n200# a_n81_n288# a_n129_n200# a_n419_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_255_n200# a_207_222# a_159_n200# a_n419_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_159_n200# a_111_n288# a_63_n200# a_n419_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n225_n200# a_n273_n288# a_n317_n200# a_n419_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X4 a_63_n200# a_15_222# a_n33_n200# a_n419_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 a_n129_n200# a_n177_222# a_n225_n200# a_n419_n374# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt diffamp_element_nodi m1_1126_642# m1_1414_418# a_890_330# m1_1318_642# m1_838_418#
+ m1_1030_418# m1_934_642# m1_1222_418# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_V6SMGN_0 m1_1030_418# a_890_330# m1_1222_418# a_890_330#
+ m1_934_642# m1_1126_642# VSUBS m1_838_418# m1_1318_642# a_890_330# a_890_330# a_890_330#
+ m1_1414_418# a_890_330# sky130_fd_pr__nfet_01v8_lvt_V6SMGN
.ends

.subckt comp_adv3 Outn bias VP OutP diffamp_element_nodi_0/a_890_330# diffamp_element_nodi_1/a_890_330#
+ VN
Xsky130_fd_pr__res_xhigh_po_2p85_8K9944_0 VP OutP VN sky130_fd_pr__res_xhigh_po_2p85_8K9944
Xsky130_fd_pr__res_xhigh_po_2p85_8K9944_1 VP Outn VN sky130_fd_pr__res_xhigh_po_2p85_8K9944
Xdiffamp_element_nodi_0 OutP m2_720_n160# diffamp_element_nodi_0/a_890_330# OutP m2_720_n160#
+ m2_720_n160# OutP m2_720_n160# VN diffamp_element_nodi
Xdiffamp_element_nodi_1 Outn m2_720_n160# diffamp_element_nodi_1/a_890_330# Outn m2_720_n160#
+ m2_720_n160# Outn m2_720_n160# VN diffamp_element_nodi
Xcurrm_comp_0 VN bias bias VN VN bias VN m2_720_n160# bias m2_720_n160# VN VN m2_720_n160#
+ bias bias bias bias m2_720_n160# bias bias VN bias VN m2_720_n160# VN bias currm_comp
.ends

.subckt sky130_fd_pr__pfet_01v8_XJ7GBL a_n33_n147# a_n73_n50# w_n211_n269# a_15_n50#
X0 a_15_n50# a_n33_n147# a_n73_n50# w_n211_n269# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_U47ZGH a_n221_n200# a_n129_n200# a_63_n200# a_15_n297#
+ a_n81_231# w_n359_n419# a_n177_n297# a_n33_n200# a_159_n200# a_111_231#
X0 a_159_n200# a_111_231# a_63_n200# w_n359_n419# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_63_n200# a_15_n297# a_n33_n200# w_n359_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_n129_n200# a_n177_n297# a_n221_n200# w_n359_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X3 a_n33_n200# a_n81_231# a_n129_n200# w_n359_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_GV8PGY a_15_n200# a_n33_222# a_111_n200# a_n81_n200#
+ a_n129_n288# a_63_n288# a_n275_n374# a_n173_n200#
X0 a_n81_n200# a_n129_n288# a_n173_n200# a_n275_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X1 a_15_n200# a_n33_222# a_n81_n200# a_n275_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X2 a_111_n200# a_63_n288# a_15_n200# a_n275_n374# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_X4XKHL a_63_n200# a_15_231# a_n33_n200# w_n263_n419#
+ a_n81_n297# a_n125_n200#
X0 a_63_n200# a_15_231# a_n33_n200# w_n263_n419# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n33_n200# a_n81_n297# a_n125_n200# w_n263_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_LH2JGW a_n81_n288# a_63_n200# a_n33_n200# a_15_222#
+ a_n227_n374# a_n125_n200#
X0 a_n33_n200# a_n81_n288# a_n125_n200# a_n227_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X1 a_63_n200# a_15_222# a_n33_n200# a_n227_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_YT8PGU a_15_n200# a_n175_n374# a_n73_n200# a_n33_n288#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n175_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PL8DH5 a_n1209_n200# a_262_n288# a_n328_n288# a_1033_n200#
+ a_n501_n200# a_n855_n200# a_616_n288# a_561_n200# a_144_n288# a_n383_n200# a_498_n288#
+ a_915_n200# a_n1154_n288# a_n737_n200# a_443_n200# a_n1311_n374# a_797_n200# a_n265_n200#
+ a_n800_n288# a_n1036_n288# a_n619_n200# a_26_n288# a_325_n200# a_n682_n288# a_679_n200#
+ a_n147_n200# a_970_n288# a_n1091_n200# a_207_n200# a_n210_n288# a_n564_n288# a_852_n288#
+ a_n918_n288# a_n29_n200# a_380_n288# a_n92_n288# a_89_n200# a_n446_n288# a_1151_n200#
+ a_734_n288# a_n973_n200# a_1088_n288#
X0 a_n29_n200# a_n92_n288# a_n147_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X1 a_915_n200# a_852_n288# a_797_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X2 a_n619_n200# a_n682_n288# a_n737_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X3 a_n855_n200# a_n918_n288# a_n973_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X4 a_325_n200# a_262_n288# a_207_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X5 a_561_n200# a_498_n288# a_443_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X6 a_n265_n200# a_n328_n288# a_n383_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X7 a_1151_n200# a_1088_n288# a_1033_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X8 a_797_n200# a_734_n288# a_679_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X9 a_89_n200# a_26_n288# a_n29_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X10 a_207_n200# a_144_n288# a_89_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X11 a_n1091_n200# a_n1154_n288# a_n1209_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=300000u
X12 a_n501_n200# a_n564_n288# a_n619_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=300000u
X13 a_n147_n200# a_n210_n288# a_n265_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X14 a_679_n200# a_616_n288# a_561_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X15 a_1033_n200# a_970_n288# a_915_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X16 a_n737_n200# a_n800_n288# a_n855_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X17 a_n973_n200# a_n1036_n288# a_n1091_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X18 a_443_n200# a_380_n288# a_325_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X19 a_n383_n200# a_n446_n288# a_n501_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
.ends

.subckt comp_to_logic Out VP In_p In_n I_Bias VSUBS
Xsky130_fd_pr__pfet_01v8_XJ7GBL_1 VM6D VM1D VP VP sky130_fd_pr__pfet_01v8_XJ7GBL
Xsky130_fd_pr__pfet_01v8_XJ7GBL_0 VM1D VP VP VM6D sky130_fd_pr__pfet_01v8_XJ7GBL
Xsky130_fd_pr__pfet_01v8_U47ZGH_0 VP VM11D VM11D VM1D VM1D VP VM1D VP VP VM1D sky130_fd_pr__pfet_01v8_U47ZGH
Xsky130_fd_pr__nfet_01v8_GV8PGY_0 VSUBS VM11D VM11D VM11D VM11D VM11D VSUBS VSUBS
+ sky130_fd_pr__nfet_01v8_GV8PGY
Xsky130_fd_pr__pfet_01v8_U47ZGH_1 VP VM12D VM12D VM6D VM6D VP VM6D VP VP VM6D sky130_fd_pr__pfet_01v8_U47ZGH
Xsky130_fd_pr__nfet_01v8_GV8PGY_1 VSUBS VM11D VM12D VM12D VM11D VM11D VSUBS VSUBS
+ sky130_fd_pr__nfet_01v8_GV8PGY
Xsky130_fd_pr__pfet_01v8_U47ZGH_2 VP VM13D VM13D VM17D VM17D VP VM17D VP VP VM17D
+ sky130_fd_pr__pfet_01v8_U47ZGH
Xsky130_fd_pr__pfet_01v8_U47ZGH_3 VP Out Out VM13D VM13D VP VM13D VP VP VM13D sky130_fd_pr__pfet_01v8_U47ZGH
Xsky130_fd_pr__pfet_01v8_X4XKHL_0 VP VM1D VM1D VP VM1D VP sky130_fd_pr__pfet_01v8_X4XKHL
Xsky130_fd_pr__pfet_01v8_X4XKHL_2 VP VM12D VM17D VP VM12D VP sky130_fd_pr__pfet_01v8_X4XKHL
Xsky130_fd_pr__pfet_01v8_X4XKHL_1 VP VM6D VM6D VP VM6D VP sky130_fd_pr__pfet_01v8_X4XKHL
Xsky130_fd_pr__nfet_01v8_lvt_LH2JGW_0 In_n VM4D VM1D In_n VSUBS VM4D sky130_fd_pr__nfet_01v8_lvt_LH2JGW
Xsky130_fd_pr__nfet_01v8_lvt_LH2JGW_2 VM13D VSUBS Out VM13D VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt_LH2JGW
Xsky130_fd_pr__nfet_01v8_lvt_LH2JGW_1 In_p VM4D VM6D In_p VSUBS VM4D sky130_fd_pr__nfet_01v8_lvt_LH2JGW
Xsky130_fd_pr__nfet_01v8_lvt_LH2JGW_3 VM17D VSUBS VM13D VM17D VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt_LH2JGW
Xsky130_fd_pr__nfet_01v8_YT8PGU_0 VM17D VSUBS VSUBS VM12D sky130_fd_pr__nfet_01v8_YT8PGU
Xsky130_fd_pr__nfet_01v8_PL8DH5_0 VSUBS I_Bias I_Bias VSUBS VM4D VSUBS I_Bias VSUBS
+ I_Bias VSUBS I_Bias VM4D VSUBS VM4D VM4D VSUBS VSUBS VM4D I_Bias I_Bias VSUBS I_Bias
+ VSUBS I_Bias VM4D VSUBS I_Bias VSUBS VM4D I_Bias I_Bias I_Bias I_Bias VM4D I_Bias
+ I_Bias VSUBS I_Bias VSUBS I_Bias I_Bias VSUBS sky130_fd_pr__nfet_01v8_PL8DH5
.ends

.subckt comparator comp_adv3_4/bias VP comp_adv3_2/bias comp_adv3_di_0/bias InRef
+ comp_to_logic_0/I_Bias comp_adv3_3/bias comp_to_logic_0/Out In VN
Xsky130_fd_pr__res_xhigh_po_0p35_Z7KPPL_0 VN m1_n2250_2600# m1_n3200_150# m1_n2870_2590#
+ m1_n2560_340# m1_n3200_150# m1_n2560_340# comp_adv3_0/OutP m1_n2870_2590# sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL
Xsky130_fd_pr__res_xhigh_po_0p35_Z7KPPL_1 VN m1_n8540_2590# m1_n9500_160# m1_n9180_2590#
+ m1_n8860_160# m1_n9500_160# m1_n8860_160# m1_n9490_2240# m1_n9180_2590# sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL
Xsky130_fd_pr__res_xhigh_po_0p35_Z7KPPL_2 VN InRef m1_n8150_160# m1_n7830_2600# m1_n7520_160#
+ m1_n8150_160# m1_n7520_160# m1_n8540_2590# m1_n7830_2600# sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL
Xcomp_adv3_di_0 comp_adv3_di_0/Outn comp_adv3_di_0/bias VP m1_n2250_2600# comp_adv3_0/OutP
+ comp_adv3_di_0/Outp VN comp_adv3_di
Xsky130_fd_pr__cap_mim_m3_2_MJMGTW_0 VN m1_n8540_2590# sky130_fd_pr__cap_mim_m3_2_MJMGTW
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0 m1_n2250_2600# comp_adv3_0/Outn sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_1 m1_n9490_2240# In sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xcomp_adv3_0 comp_adv3_0/Outn comp_adv3_0/bias VP comp_adv3_0/OutP comp_adv3_1/OutP
+ comp_adv3_1/Outn VN comp_adv3
Xcomp_adv3_1 comp_adv3_1/Outn comp_adv3_1/bias VP comp_adv3_1/OutP m1_n8540_2590#
+ m1_n9490_2240# VN comp_adv3
Xcomp_adv3_2 comp_adv3_2/Outn comp_adv3_2/bias VP comp_adv3_2/OutP comp_adv3_di_0/Outp
+ comp_adv3_di_0/Outn VN comp_adv3
Xcomp_to_logic_0 comp_to_logic_0/Out VP comp_adv3_4/OutP comp_adv3_4/Outn comp_to_logic_0/I_Bias
+ VN comp_to_logic
Xcomp_adv3_3 comp_adv3_3/Outn comp_adv3_3/bias VP comp_adv3_3/OutP comp_adv3_2/OutP
+ comp_adv3_2/Outn VN comp_adv3
Xcomp_adv3_4 comp_adv3_4/Outn comp_adv3_4/bias VP comp_adv3_4/OutP comp_adv3_3/OutP
+ comp_adv3_3/Outn VN comp_adv3
.ends

.subckt sky130_fd_pr__nfet_01v8_PJG2KG a_50_n200# a_n108_n200# a_n50_n288# a_n210_n374#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n210_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_82JNGJ a_n221_n200# a_n129_n200# a_63_n200# a_111_222#
+ a_n33_n200# a_15_n288# a_n81_222# a_n177_n288# a_159_n200# a_n323_n374#
X0 a_n33_n200# a_n81_222# a_n129_n200# a_n323_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_159_n200# a_111_222# a_63_n200# a_n323_n374# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_63_n200# a_15_n288# a_n33_n200# a_n323_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 a_n129_n200# a_n177_n288# a_n221_n200# a_n323_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
.ends

.subckt currm_n m1_68_150# m1_164_390# a_122_62# VSUBS
Xsky130_fd_pr__nfet_01v8_PJG2KG_0 VSUBS m1_68_150# a_122_62# VSUBS sky130_fd_pr__nfet_01v8_PJG2KG
Xsky130_fd_pr__nfet_01v8_82JNGJ_0 m1_68_150# m1_164_390# m1_164_390# a_122_62# m1_68_150#
+ a_122_62# a_122_62# a_122_62# m1_68_150# VSUBS sky130_fd_pr__nfet_01v8_82JNGJ
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4LMUGG a_355_n200# a_413_n297# a_n285_n200# a_29_n297#
+ a_n227_n297# a_285_n297# a_227_n200# a_n157_n200# a_n541_n200# w_n679_n419# a_n483_n297#
+ a_n99_n297# a_483_n200# a_157_n297# a_99_n200# a_n413_n200# a_n29_n200# a_n355_n297#
X0 a_227_n200# a_157_n297# a_99_n200# w_n679_n419# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=350000u
X1 a_n285_n200# a_n355_n297# a_n413_n200# w_n679_n419# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=350000u
X2 a_99_n200# a_29_n297# a_n29_n200# w_n679_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=350000u
X3 a_355_n200# a_285_n297# a_227_n200# w_n679_n419# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=350000u
X4 a_483_n200# a_413_n297# a_355_n200# w_n679_n419# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=350000u
X5 a_n29_n200# a_n99_n297# a_n157_n200# w_n679_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=350000u
X6 a_n413_n200# a_n483_n297# a_n541_n200# w_n679_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=350000u
X7 a_n157_n200# a_n227_n297# a_n285_n200# w_n679_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_LKHJAY a_29_n297# a_n287_n200# a_n229_n297# a_229_n200#
+ w_n425_n419# a_n29_n200#
X0 a_229_n200# a_29_n297# a_n29_n200# w_n425_n419# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X1 a_n29_n200# a_n229_n297# a_n287_n200# w_n425_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
.ends

.subckt currm_p m1_60_n360# m1_70_460# m1_190_n590# m1_n50_n680#
Xsky130_fd_pr__pfet_01v8_lvt_4LMUGG_0 m1_190_n590# m1_n50_n680# m1_60_n360# m1_n50_n680#
+ m1_n50_n680# m1_n50_n680# m1_60_n360# m1_190_n590# m1_60_n360# m1_70_460# m1_n50_n680#
+ m1_n50_n680# m1_60_n360# m1_n50_n680# m1_190_n590# m1_190_n590# m1_60_n360# m1_n50_n680#
+ sky130_fd_pr__pfet_01v8_lvt_4LMUGG
Xsky130_fd_pr__pfet_01v8_lvt_LKHJAY_0 m1_n50_n680# m1_70_460# m1_n50_n680# m1_70_460#
+ m1_70_460# m1_60_n360# sky130_fd_pr__pfet_01v8_lvt_LKHJAY
.ends

.subckt sky130_fd_pr__pfet_01v8_PD4XN5 a_29_n297# a_n129_n297# a_129_n200# w_n325_n419#
+ a_n29_n200# a_n187_n200#
X0 a_129_n200# a_29_n297# a_n29_n200# w_n325_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_n29_n200# a_n129_n297# a_n187_n200# w_n325_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_U4PWGH a_n129_n200# a_63_n200# a_n225_n200# a_15_n297#
+ a_n81_231# a_n177_n297# a_n273_231# a_n321_n200# w_n551_n419# a_n33_n200# a_159_n200#
+ a_n413_n200# a_111_231# a_255_n200# a_207_n297# a_351_n200# a_n369_n297# a_303_231#
X0 a_255_n200# a_207_n297# a_159_n200# w_n551_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n321_n200# a_n369_n297# a_n413_n200# w_n551_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X2 a_159_n200# a_111_231# a_63_n200# w_n551_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n225_n200# a_n273_231# a_n321_n200# w_n551_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X4 a_63_n200# a_15_n297# a_n33_n200# w_n551_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_n129_n200# a_n177_n297# a_n225_n200# w_n551_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X6 a_351_n200# a_303_231# a_255_n200# w_n551_n419# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X7 a_n33_n200# a_n81_231# a_n129_n200# w_n551_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt currm_ps m1_170_170# a_132_72# w_132_72# m1_80_400#
Xsky130_fd_pr__pfet_01v8_PD4XN5_0 a_132_72# a_132_72# w_132_72# w_132_72# m1_80_400#
+ w_132_72# sky130_fd_pr__pfet_01v8_PD4XN5
Xsky130_fd_pr__pfet_01v8_U4PWGH_0 m1_170_170# m1_170_170# m1_80_400# a_132_72# a_132_72#
+ a_132_72# a_132_72# m1_170_170# w_132_72# m1_80_400# m1_80_400# m1_80_400# a_132_72#
+ m1_170_170# a_132_72# m1_80_400# a_132_72# a_132_72# sky130_fd_pr__pfet_01v8_U4PWGH
.ends

.subckt sky130_fd_pr__nfet_01v8_6H2JYD a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_N3PKNJ c2_n3251_n1000# m4_n3351_n1100#
X0 c2_n3251_n1000# m4_n3351_n1100# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_9A2JGL a_n81_109# a_15_109# a_n225_n597# a_15_n509#
+ a_n177_n509# a_111_n509# a_207_109# a_63_n87# a_159_531# a_n371_n683# a_n33_n597#
+ a_n33_531# a_n129_n87# a_n177_109# a_n225_531# a_n81_n509# a_111_109# a_n129_21#
+ a_159_n597# a_63_21# a_n269_n509# a_n269_109# a_207_n509#
X0 a_15_109# a_n33_531# a_n81_109# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_111_109# a_63_21# a_15_109# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X2 a_n81_109# a_n129_21# a_n177_109# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n177_109# a_n225_531# a_n269_109# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X4 a_n81_n509# a_n129_n87# a_n177_n509# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_15_n509# a_n33_n597# a_n81_n509# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X6 a_207_109# a_159_531# a_111_109# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X7 a_207_n509# a_159_n597# a_111_n509# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X8 a_n177_n509# a_n225_n597# a_n269_n509# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X9 a_111_n509# a_63_n87# a_15_n509# a_n371_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_VCBWSW a_n513_n200# a_n989_n200# a_n129_n200# a_63_n200#
+ a_n225_n200# a_15_n297# a_n561_n297# a_n81_231# a_927_n200# a_n177_n297# a_879_231#
+ a_n273_231# a_n321_n200# a_639_n200# a_735_n200# a_n33_n200# a_n465_231# a_n897_n200#
+ a_831_n200# a_447_n200# a_783_n297# a_399_n297# a_543_n200# a_159_n200# a_n609_n200#
+ a_n945_n297# a_n657_231# a_495_231# a_111_231# a_255_n200# a_n705_n200# a_591_n297#
+ a_207_n297# a_351_n200# a_n801_n200# a_n849_231# a_n417_n200# a_n369_n297# a_n753_n297#
+ w_n1127_n419# a_687_231# a_303_231#
X0 a_n609_n200# a_n657_231# a_n705_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_927_n200# a_879_231# a_831_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_n897_n200# a_n945_n297# a_n989_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X3 a_255_n200# a_207_n297# a_159_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n321_n200# a_n369_n297# a_n417_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_543_n200# a_495_231# a_447_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_831_n200# a_783_n297# a_735_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_159_n200# a_111_231# a_63_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X8 a_n225_n200# a_n273_231# a_n321_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X9 a_447_n200# a_399_n297# a_351_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_n513_n200# a_n561_n297# a_n609_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_63_n200# a_15_n297# a_n33_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_735_n200# a_687_231# a_639_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X13 a_n801_n200# a_n849_231# a_n897_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X14 a_n129_n200# a_n177_n297# a_n225_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X15 a_n417_n200# a_n465_231# a_n513_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 a_639_n200# a_591_n297# a_543_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 a_n705_n200# a_n753_n297# a_n801_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 a_351_n200# a_303_231# a_255_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 a_n33_n200# a_n81_231# a_n129_n200# w_n1127_n419# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_MJMGTW#0 c2_n3251_n2000# m4_n3351_n2100#
X0 c2_n3251_n2000# m4_n3351_n2100# sky130_fd_pr__cap_mim_m3_2 l=2e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_E6B2KN a_129_n200# a_29_n288# a_n129_n288# a_n289_n374#
+ a_n29_n200# a_n187_n200#
X0 a_129_n200# a_29_n288# a_n29_n200# a_n289_n374# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_n29_n200# a_n129_n288# a_n187_n200# a_n289_n374# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_UAQRRG a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_LH2JGW#0 a_n81_n288# a_63_n200# a_n33_n200# a_15_222#
+ a_n227_n374# a_n125_n200#
X0 a_n33_n200# a_n81_n288# a_n125_n200# a_n227_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X1 a_63_n200# a_15_222# a_n33_n200# a_n227_n374# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG#4 m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt fb_dark_current VP InP InN VN
Xcurrm_n_2 m2_250_740# m1_950_1560# I_Bias VN currm_n
Xcurrm_p_5 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
Xcurrm_n_3 m2_250_740# m1_950_1560# I_Bias VN currm_n
Xcurrm_p_6 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
Xcurrm_ps_0 m1_9810_5770# m1_9810_5770# VP currm_ps_0/m1_80_400# currm_ps
Xcurrm_n_4 currm_n_4/m1_68_150# m1_n5100_670# m1_n5100_670# VN currm_n
Xcurrm_p_7 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
Xcurrm_ps_1 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_n_5 currm_n_5/m1_68_150# m1_4960_670# m1_4960_670# VN currm_n
Xsky130_fd_pr__nfet_01v8_6H2JYD_0 m1_n830_1270# Disable_FB VN VN sky130_fd_pr__nfet_01v8_6H2JYD
Xcurrm_p_9 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
Xcurrm_p_8 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
Xcurrm_ps_19 m1_n6550_3300# m1_n6550_3300# VP currm_ps_19/m1_80_400# currm_ps
Xcurrm_ps_18 m1_9390_670# m1_n6550_3300# VP currm_ps_18/m1_80_400# currm_ps
Xcurrm_ps_2 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_n_7 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xcurrm_n_6 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xcurrm_ps_3 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_n_8 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xcurrm_ps_4 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_n_9 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xcurrm_ps_5 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_p_20 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xcurrm_p_21 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xcurrm_p_10 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
Xcurrm_ps_6 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_p_11 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
Xcurrm_ps_7 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_ps_8 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_p_12 currm_p_12/m1_60_n360# VP m1_n5100_670# m1_7940_2770# currm_p
Xcurrm_p_13 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xcurrm_ps_9 Out m1_9810_5770# VP m2_9370_4730# currm_ps
Xcurrm_p_14 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xcurrm_p_15 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xcurrm_p_16 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xcurrm_p_17 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xsky130_fd_pr__cap_mim_m3_2_N3PKNJ_0 VN I_Bias sky130_fd_pr__cap_mim_m3_2_N3PKNJ
Xsky130_fd_pr__nfet_01v8_9A2JGL_1 m1_9390_670# VN Disable_FB m1_9390_670# m1_9390_670#
+ VN VN Disable_FB Disable_FB VN Disable_FB Disable_FB Disable_FB VN Disable_FB VN
+ m1_9390_670# Disable_FB Disable_FB Disable_FB VN m1_9390_670# m1_9390_670# sky130_fd_pr__nfet_01v8_9A2JGL
Xsky130_fd_pr__cap_mim_m3_2_N3PKNJ_1 VN I_Bias sky130_fd_pr__cap_mim_m3_2_N3PKNJ
Xcurrm_n_40 m2_9090_740# Out m1_9390_670# VN currm_n
Xcurrm_p_18 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xcurrm_p_19 m2_4260_3100# VP m1_9810_5770# m1_7940_2770# currm_p
Xsky130_fd_pr__pfet_01v8_VCBWSW_0 VP m1_9810_5770# VP VP m1_9810_5770# m1_n830_1270#
+ m1_n830_1270# m1_n830_1270# m1_9810_5770# m1_n830_1270# m1_n830_1270# m1_n830_1270#
+ VP VP m1_9810_5770# m1_9810_5770# m1_n830_1270# VP VP VP m1_n830_1270# m1_n830_1270#
+ m1_9810_5770# m1_9810_5770# m1_9810_5770# m1_n830_1270# m1_n830_1270# m1_n830_1270#
+ m1_n830_1270# VP VP m1_n830_1270# m1_n830_1270# m1_9810_5770# m1_9810_5770# m1_n830_1270#
+ m1_9810_5770# m1_n830_1270# m1_n830_1270# VP m1_n830_1270# m1_n830_1270# sky130_fd_pr__pfet_01v8_VCBWSW
Xcurrm_n_41 m2_9090_740# Out m1_9390_670# VN currm_n
Xsky130_fd_pr__cap_mim_m3_2_MJMGTW_0 VP VN sky130_fd_pr__cap_mim_m3_2_MJMGTW#0
Xcurrm_n_42 m2_9090_740# Out m1_9390_670# VN currm_n
Xcurrm_n_31 m2_n6460_740# m1_9390_670# m1_9390_670# VN currm_n
Xcurrm_n_20 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_n_43 currm_n_43/m1_68_150# m1_9810_5770# I_Bias VN currm_n
Xcurrm_n_10 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xcurrm_n_32 m2_9090_740# Out m1_9390_670# VN currm_n
Xcurrm_n_21 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_n_11 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xcurrm_n_12 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xcurrm_n_45 m2_200_n880# I_Bias I_Bias VN currm_n
Xcurrm_n_44 m2_200_n880# I_Bias I_Bias VN currm_n
Xcurrm_n_33 currm_n_33/m1_68_150# m1_n6550_3300# I_Bias VN currm_n
Xcurrm_n_23 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_n_22 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_n_35 m2_9090_740# Out m1_9390_670# VN currm_n
Xcurrm_n_13 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xcurrm_n_46 m2_200_n880# I_Bias I_Bias VN currm_n
Xcurrm_n_36 m2_9090_740# Out m1_9390_670# VN currm_n
Xcurrm_n_14 m2_4080_740# m1_9810_5770# m1_4960_670# VN currm_n
Xsky130_fd_pr__nfet_01v8_E6B2KN_0 m1_950_1560# InP InP VN m1_970_2720# m1_950_1560#
+ sky130_fd_pr__nfet_01v8_E6B2KN
Xcurrm_n_47 m2_200_n880# I_Bias I_Bias VN currm_n
Xsky130_fd_pr__pfet_01v8_UAQRRG_0 m1_n830_1270# VP VP Disable_FB sky130_fd_pr__pfet_01v8_UAQRRG
Xcurrm_n_37 m2_9090_740# Out m1_9390_670# VN currm_n
Xsky130_fd_pr__nfet_01v8_E6B2KN_1 m1_950_1560# InN InN VN m1_7940_2770# m1_950_1560#
+ sky130_fd_pr__nfet_01v8_E6B2KN
Xsky130_fd_pr__nfet_01v8_lvt_LH2JGW_0 Disable_FB VN I_Bias Disable_FB VN VN sky130_fd_pr__nfet_01v8_lvt_LH2JGW#0
Xcurrm_n_15 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_n_38 m2_9090_740# Out m1_9390_670# VN currm_n
Xcurrm_n_16 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_n_39 m2_9090_740# Out m1_9390_670# VN currm_n
Xcurrm_n_17 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_n_18 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_n_19 m2_n5090_n880# m1_n6550_3300# m1_n5100_670# VN currm_n
Xcurrm_p_0 currm_p_0/m1_60_n360# VP m1_970_2720# m1_970_2720# currm_p
Xcurrm_p_1 currm_p_1/m1_60_n360# VP m1_7940_2770# m1_7940_2770# currm_p
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_2 m1_970_2720# VP sky130_fd_pr__cap_mim_m3_2_LJ5JLG#4
Xcurrm_p_2 currm_p_2/m1_60_n360# VP m1_4960_670# m1_970_2720# currm_p
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_3 m1_7940_2770# VP sky130_fd_pr__cap_mim_m3_2_LJ5JLG#4
Xcurrm_n_0 m2_250_740# m1_950_1560# I_Bias VN currm_n
Xcurrm_p_3 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
Xcurrm_n_1 m2_250_740# m1_950_1560# I_Bias VN currm_n
Xcurrm_p_4 m2_n5120_4740# VP m1_n6550_3300# m1_970_2720# currm_p
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WXTTNJ#0 c1_n2050_n2000# m3_n2150_n2100#
X0 c1_n2050_n2000# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_834VMG a_2487_n400# a_n29_n400# a_n2487_n488# a_1229_n400#
+ a_n2647_n574# a_n2545_n400# a_n1229_n488# a_1287_n488# a_n1287_n400# a_29_n488#
X0 a_n29_n400# a_n1229_n488# a_n1287_n400# a_n2647_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X1 a_n1287_n400# a_n2487_n488# a_n2545_n400# a_n2647_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X2 a_1229_n400# a_29_n488# a_n29_n400# a_n2647_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
X3 a_2487_n400# a_1287_n488# a_1229_n400# a_n2647_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_26RGPZ a_n225_n909# a_n129_109# a_n369_21# a_n465_931#
+ a_447_109# a_399_21# a_n321_n909# a_n177_n87# a_n81_n997# a_n321_109# a_n509_109#
+ a_n33_n909# a_n509_n909# a_159_109# a_n369_n87# a_111_931# a_447_n909# a_351_109#
+ a_n33_109# a_n611_n1083# a_159_n909# a_303_n997# a_n225_109# a_303_931# a_n177_21#
+ a_255_n909# a_399_n87# a_n465_n997# a_207_21# a_351_n909# a_n417_n909# a_63_109#
+ a_n81_931# a_15_n87# a_15_21# a_111_n997# a_n417_109# a_n273_931# a_n129_n909# a_n273_n997#
+ a_255_109# a_207_n87# a_63_n909#
X0 a_351_n909# a_303_n997# a_255_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X1 a_n33_n909# a_n81_n997# a_n129_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X2 a_255_n909# a_207_n87# a_159_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X3 a_n33_109# a_n81_931# a_n129_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X4 a_n321_n909# a_n369_n87# a_n417_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X5 a_351_109# a_303_931# a_255_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X6 a_159_109# a_111_931# a_63_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X7 a_255_109# a_207_21# a_159_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8 a_447_109# a_399_21# a_351_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.24e+12p pd=8.62e+06u as=0p ps=0u w=4e+06u l=150000u
X9 a_n321_109# a_n369_21# a_n417_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X10 a_n417_109# a_n465_931# a_n509_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.24e+12p ps=8.62e+06u w=4e+06u l=150000u
X11 a_n225_109# a_n273_931# a_n321_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=0p ps=0u w=4e+06u l=150000u
X12 a_n129_109# a_n177_21# a_n225_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 a_159_n909# a_111_n997# a_63_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.32e+12p ps=8.66e+06u w=4e+06u l=150000u
X14 a_n225_n909# a_n273_n997# a_n321_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=8.66e+06u as=0p ps=0u w=4e+06u l=150000u
X15 a_447_n909# a_399_n87# a_351_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.24e+12p pd=8.62e+06u as=0p ps=0u w=4e+06u l=150000u
X16 a_63_n909# a_15_n87# a_n33_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X17 a_63_109# a_15_21# a_n33_109# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 a_n129_n909# a_n177_n87# a_n225_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 a_n417_n909# a_n465_n997# a_n509_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.24e+12p ps=8.62e+06u w=4e+06u l=150000u
.ends

.subckt isource_conv_tsmal m1_4500_6730# m1_4590_7330# m1_4410_6620# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_26RGPZ_0 m1_4590_7330# m1_4500_6730# m1_4410_6620# m1_4410_6620#
+ m1_4500_6730# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4410_6620# m1_4500_6730#
+ m1_4500_6730# m1_4590_7330# m1_4500_6730# m1_4590_7330# m1_4410_6620# m1_4410_6620#
+ m1_4500_6730# m1_4590_7330# m1_4590_7330# VSUBS m1_4590_7330# m1_4410_6620# m1_4590_7330#
+ m1_4410_6620# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4410_6620# m1_4410_6620#
+ m1_4590_7330# m1_4590_7330# m1_4500_6730# m1_4410_6620# m1_4410_6620# m1_4410_6620#
+ m1_4410_6620# m1_4590_7330# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4500_6730#
+ m1_4410_6620# m1_4500_6730# sky130_fd_pr__nfet_01v8_lvt_26RGPZ
.ends

.subckt sky130_fd_pr__nfet_01v8_HZ8P49 a_2487_n400# a_n6261_n488# a_n29_n400# a_5003_n400#
+ a_3803_n488# a_n2487_n488# a_n3803_n400# a_n6421_n574# a_1229_n400# a_n5003_n488#
+ a_2545_n488# a_n2545_n400# a_n1229_n488# a_5061_n488# a_n5061_n400# a_3745_n400#
+ a_1287_n488# a_6261_n400# a_n1287_n400# a_29_n488# a_n6319_n400# a_n3745_n488#
X0 a_6261_n400# a_5061_n488# a_5003_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X1 a_n29_n400# a_n1229_n488# a_n1287_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X2 a_n2545_n400# a_n3745_n488# a_n3803_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X3 a_n1287_n400# a_n2487_n488# a_n2545_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4 a_5003_n400# a_3803_n488# a_3745_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X5 a_n3803_n400# a_n5003_n488# a_n5061_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X6 a_1229_n400# a_29_n488# a_n29_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
X7 a_3745_n400# a_2545_n488# a_2487_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X8 a_n5061_n400# a_n6261_n488# a_n6319_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X9 a_2487_n400# a_1287_n488# a_1229_n400# a_n6421_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
.ends

.subckt isource_ref_transistor m1_n370_110# m1_887_21# m1_890_680# VSUBS
Xsky130_fd_pr__nfet_01v8_HZ8P49_0 m1_890_680# m1_887_21# m1_890_680# m1_890_680# m1_887_21#
+ m1_887_21# m1_n370_110# VSUBS m1_n370_110# m1_887_21# m1_887_21# m1_890_680# m1_887_21#
+ m1_887_21# m1_890_680# m1_n370_110# m1_887_21# m1_n370_110# m1_n370_110# m1_887_21#
+ m1_n370_110# m1_887_21# sky130_fd_pr__nfet_01v8_HZ8P49
.ends

.subckt sky130_fd_pr__pfet_01v8_ACY9XJ#0#0 a_20_n918# a_20_118# a_n78_n918# a_n33_21#
+ a_n78_118# w_n216_n1137# a_n33_n1015#
X0 a_20_118# a_n33_21# a_n78_118# w_n216_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X1 a_20_n918# a_n33_n1015# a_n78_n918# w_n216_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
.ends

.subckt sky130_fd_pr__pfet_01v8_J24RLQ#0#0 a_n416_118# a_n100_n1015# a_358_118# a_n416_n918#
+ a_n674_118# a_n158_118# a_n100_21# a_158_n1015# a_n358_21# w_n812_n1137# a_158_21#
+ a_358_n918# a_416_n1015# a_n358_n1015# a_100_n918# a_n674_n918# a_n616_21# a_416_21#
+ a_n616_n1015# a_n158_n918# a_616_118# a_100_118# a_616_n918#
X0 a_100_118# a_n100_21# a_n158_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X1 a_616_n918# a_416_n1015# a_358_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X2 a_358_n918# a_158_n1015# a_100_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X3 a_616_118# a_416_21# a_358_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X4 a_100_n918# a_n100_n1015# a_n158_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X5 a_358_118# a_158_21# a_100_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 a_n416_118# a_n616_21# a_n674_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X7 a_n416_n918# a_n616_n1015# a_n674_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X8 a_n158_n918# a_n358_n1015# a_n416_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 a_n158_118# a_n358_21# a_n416_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
.ends

.subckt isource_cmirror#0 m1_0_1060# li_0_0# m1_110_820#
Xsky130_fd_pr__pfet_01v8_ACY9XJ_0 m1_250_820# m1_250_820# m1_110_820# m1_0_1060# m1_110_820#
+ li_0_0# m1_0_1060# sky130_fd_pr__pfet_01v8_ACY9XJ#0#0
Xsky130_fd_pr__pfet_01v8_J24RLQ_0 li_0_0# m1_0_1060# m1_250_820# li_0_0# m1_250_820#
+ m1_250_820# m1_0_1060# m1_0_1060# m1_0_1060# li_0_0# m1_0_1060# m1_250_820# m1_0_1060#
+ m1_0_1060# li_0_0# m1_250_820# m1_0_1060# m1_0_1060# m1_0_1060# m1_250_820# li_0_0#
+ li_0_0# li_0_0# sky130_fd_pr__pfet_01v8_J24RLQ#0#0
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_JAGHGM a_n1331_n1562# a_n671_1000# a_919_n1432#
+ a_389_n1432# a_n141_1000# a_919_1000# a_389_1000# a_n141_n1432# a_n1201_n1432# a_n1201_1000#
+ a_n671_n1432#
X0 a_n1201_n1432# a_n1201_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1 a_919_n1432# a_919_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X2 a_n671_n1432# a_n671_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3 a_n141_n1432# a_n141_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X4 a_389_n1432# a_389_1000# a_n1331_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
.ends

.subckt isource_out m1_18730_12160# isource_cmirror_0/m1_0_1060# m1_21256_12488# m1_20970_12680#
+ li_23190_12600# VSUBS isource_conv_tsmal_0/m1_4500_6730#
Xsky130_fd_pr__nfet_01v8_834VMG_0 VSUBS VSUBS m1_21256_12488# m1_18730_12160# VSUBS
+ VSUBS m1_21256_12488# m1_21256_12488# m1_18730_12160# m1_21256_12488# sky130_fd_pr__nfet_01v8_834VMG
Xisource_conv_tsmal_0 isource_conv_tsmal_0/m1_4500_6730# m1_16760_11560# m1_20970_12680#
+ VSUBS isource_conv_tsmal
Xisource_ref_transistor_0 m1_18730_12160# m1_16760_11560# m1_20970_12680# VSUBS isource_ref_transistor
Xisource_cmirror_0 isource_cmirror_0/m1_0_1060# li_23190_12600# m1_20970_12680# isource_cmirror#0
Xisource_ref_transistor_1 m1_20970_12680# m1_16760_11560# m1_18730_12160# VSUBS isource_ref_transistor
Xsky130_fd_pr__res_xhigh_po_1p41_JAGHGM_0 VSUBS m1_23460_11560# VSUBS m1_24000_9140#
+ m1_23460_11560# m1_24520_11560# m1_24520_11560# m1_24000_9140# m1_22920_9140# m1_16760_11560#
+ m1_22920_9140# sky130_fd_pr__res_xhigh_po_1p41_JAGHGM
.ends

.subckt isource_conv_tsmal_nwell m1_4500_6730# m1_4590_7330# w_4356_6496# dw_4150_6290#
+ m1_4410_6620#
Xsky130_fd_pr__nfet_01v8_lvt_26RGPZ_0 m1_4590_7330# m1_4500_6730# m1_4410_6620# m1_4410_6620#
+ m1_4500_6730# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4410_6620# m1_4500_6730#
+ m1_4500_6730# m1_4590_7330# m1_4500_6730# m1_4590_7330# m1_4410_6620# m1_4410_6620#
+ m1_4500_6730# m1_4590_7330# m1_4590_7330# w_4356_6496# m1_4590_7330# m1_4410_6620#
+ m1_4590_7330# m1_4410_6620# m1_4410_6620# m1_4500_6730# m1_4410_6620# m1_4410_6620#
+ m1_4410_6620# m1_4590_7330# m1_4590_7330# m1_4500_6730# m1_4410_6620# m1_4410_6620#
+ m1_4410_6620# m1_4410_6620# m1_4590_7330# m1_4410_6620# m1_4500_6730# m1_4410_6620#
+ m1_4500_6730# m1_4410_6620# m1_4500_6730# sky130_fd_pr__nfet_01v8_lvt_26RGPZ
.ends

.subckt sky130_fd_pr__pfet_01v8_QDYTZD a_n200_n147# a_n258_n50# w_n396_n269# a_200_n50#
X0 a_200_n50# a_n200_n147# a_n258_n50# w_n396_n269# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_U3V43Z a_n258_n50# a_n200_n138# a_n360_n224# a_200_n50#
X0 a_200_n50# a_n200_n138# a_n258_n50# a_n360_n224# sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_E9U3PA a_363_n400# a_114_n488# a_n29_n400# a_408_422#
+ a_n278_n488# a_461_n400# a_n127_n400# a_n180_422# a_n82_n488# a_16_422# a_n225_n400#
+ a_310_n488# a_n519_n400# a_69_n400# a_n323_n400# a_n474_n488# a_212_422# a_167_n400#
+ a_n376_422# a_n421_n400# a_265_n400# a_n621_n574#
X0 a_n421_n400# a_n474_n488# a_n519_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X1 a_461_n400# a_408_422# a_363_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X2 a_n127_n400# a_n180_422# a_n225_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X3 a_167_n400# a_114_n488# a_69_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X4 a_n225_n400# a_n278_n488# a_n323_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X5 a_265_n400# a_212_422# a_167_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=200000u
X6 a_69_n400# a_16_422# a_n29_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X7 a_n323_n400# a_n376_422# a_n421_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X8 a_n29_n400# a_n82_n488# a_n127_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X9 a_363_n400# a_310_n488# a_265_n400# a_n621_n574# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
.ends

.subckt isource_startup li_2190_920# m1_360_100# sky130_fd_pr__nfet_01v8_U3V43Z_0/a_200_n50#
+ VSUBS
Xsky130_fd_pr__pfet_01v8_QDYTZD_1 m1_360_100# m1_330_800# li_2190_920# li_2190_920#
+ sky130_fd_pr__pfet_01v8_QDYTZD
Xsky130_fd_pr__nfet_01v8_U3V43Z_0 VSUBS m1_330_800# VSUBS sky130_fd_pr__nfet_01v8_U3V43Z_0/a_200_n50#
+ sky130_fd_pr__nfet_01v8_U3V43Z
Xsky130_fd_pr__nfet_01v8_lvt_E9U3PA_0 VSUBS m1_360_100# VSUBS m1_360_100# m1_360_100#
+ m1_330_800# m1_330_800# m1_360_100# m1_360_100# m1_360_100# VSUBS m1_360_100# m1_330_800#
+ m1_330_800# m1_330_800# m1_360_100# m1_360_100# VSUBS m1_360_100# VSUBS m1_330_800#
+ VSUBS sky130_fd_pr__nfet_01v8_lvt_E9U3PA
.ends

.subckt isource_ref_5transistors m2_12120_850# m1_12450_1060# m2_220_270# VSUBS
Xisource_ref_transistor_0 m2_220_270# m1_12450_1060# m2_12120_850# VSUBS isource_ref_transistor
Xisource_ref_transistor_1 VSUBS m1_12450_1060# m1_12450_1060# VSUBS isource_ref_transistor
Xisource_ref_transistor_3 m2_220_270# m1_12450_1060# m2_12120_850# VSUBS isource_ref_transistor
Xisource_ref_transistor_4 m2_220_270# m1_12450_1060# m2_12120_850# VSUBS isource_ref_transistor
.ends

.subckt sky130_fd_pr__nfet_01v8_TV3VM6 a_n658_n400# a_n3276_n574# a_n600_n488# a_n3174_n400#
+ a_1858_n400# a_n1858_n488# a_3116_n400# a_1916_n488# a_658_n488# a_600_n400# a_n1916_n400#
+ a_n3116_n488#
X0 a_1858_n400# a_658_n488# a_600_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X1 a_n658_n400# a_n1858_n488# a_n1916_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X2 a_n1916_n400# a_n3116_n488# a_n3174_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X3 a_3116_n400# a_1916_n488# a_1858_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
X4 a_600_n400# a_n600_n488# a_n658_n400# a_n3276_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_WY4VMC a_n29_n400# a_1229_n400# a_n1229_n488# a_n1389_n574#
+ a_n1287_n400# a_29_n488#
X0 a_n29_n400# a_n1229_n488# a_n1287_n400# a_n1389_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=6e+06u
X1 a_1229_n400# a_29_n488# a_n29_n400# a_n1389_n574# sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=6e+06u
.ends

.subckt isource_ref m2_12700_7520# m1_1370_6840# m1_12708_6228# m1_5600_140# m1_130_6460#
+ VSUBS
Xisource_ref_transistor_0 VSUBS m1_5600_140# m1_5600_140# VSUBS isource_ref_transistor
Xisource_ref_5transistors_0 m1_1370_6840# m1_5600_140# m1_130_6460# VSUBS isource_ref_5transistors
Xisource_ref_5transistors_1 m1_1370_6840# m1_5600_140# m1_130_6460# VSUBS isource_ref_5transistors
Xsky130_fd_pr__nfet_01v8_TV3VM6_0 m1_130_6460# VSUBS m1_5600_140# m1_130_6460# m1_130_6460#
+ m1_5600_140# m1_1370_6840# m1_5600_140# m1_5600_140# m1_1370_6840# m1_1370_6840#
+ m1_5600_140# sky130_fd_pr__nfet_01v8_TV3VM6
Xsky130_fd_pr__nfet_01v8_WY4VMC_0 m1_130_6460# VSUBS m1_12708_6228# VSUBS VSUBS m1_12708_6228#
+ sky130_fd_pr__nfet_01v8_WY4VMC
.ends

.subckt sky130_fd_pr__pfet_01v8_ACY9XJ#0 a_20_n918# a_20_118# a_n78_n918# a_n33_21#
+ a_n78_118# w_n216_n1137# a_n33_n1015#
X0 a_20_118# a_n33_21# a_n78_118# w_n216_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
X1 a_20_n918# a_n33_n1015# a_n78_n918# w_n216_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=200000u
.ends

.subckt sky130_fd_pr__pfet_01v8_J24RLQ#0 a_n416_118# a_n100_n1015# a_358_118# a_n416_n918#
+ a_n674_118# a_n158_118# a_n100_21# a_158_n1015# a_n358_21# w_n812_n1137# a_158_21#
+ a_358_n918# a_416_n1015# a_n358_n1015# a_100_n918# a_n674_n918# a_n616_21# a_416_21#
+ a_n616_n1015# a_n158_n918# a_616_118# a_100_118# a_616_n918#
X0 a_100_118# a_n100_21# a_n158_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X1 a_616_n918# a_416_n1015# a_358_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X2 a_358_n918# a_158_n1015# a_100_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X3 a_616_118# a_416_21# a_358_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X4 a_100_n918# a_n100_n1015# a_n158_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X5 a_358_118# a_158_21# a_100_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 a_n416_118# a_n616_21# a_n674_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X7 a_n416_n918# a_n616_n1015# a_n674_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X8 a_n158_n918# a_n358_n1015# a_n416_n918# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 a_n158_118# a_n358_21# a_n416_118# w_n812_n1137# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
.ends

.subckt isource_cmirror m1_0_1060# li_0_0# m1_250_820# m1_110_820#
Xsky130_fd_pr__pfet_01v8_ACY9XJ_0 m1_250_820# m1_250_820# m1_110_820# m1_0_1060# m1_110_820#
+ li_0_0# m1_0_1060# sky130_fd_pr__pfet_01v8_ACY9XJ#0
Xsky130_fd_pr__pfet_01v8_J24RLQ_0 li_0_0# m1_0_1060# m1_250_820# li_0_0# m1_250_820#
+ m1_250_820# m1_0_1060# m1_0_1060# m1_0_1060# li_0_0# m1_0_1060# m1_250_820# m1_0_1060#
+ m1_0_1060# li_0_0# m1_250_820# m1_0_1060# m1_0_1060# m1_0_1060# m1_250_820# li_0_0#
+ li_0_0# li_0_0# sky130_fd_pr__pfet_01v8_J24RLQ#0
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_BQY2W7 a_n406_1000# a_n1996_1000# a_n1996_n1432#
+ a_654_n1432# a_1714_1000# a_1714_n1432# a_1184_n1432# a_n1466_1000# a_1184_1000#
+ a_n2126_n1562# a_n406_n1432# a_654_1000# a_n936_1000# a_n936_n1432# a_n1466_n1432#
+ a_124_n1432# a_124_1000#
X0 a_654_n1432# a_654_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1 a_124_n1432# a_124_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X2 a_n1996_n1432# a_n1996_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X3 a_n1466_n1432# a_n1466_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X4 a_n936_n1432# a_n936_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X5 a_1714_n1432# a_1714_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X6 a_n406_n1432# a_n406_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X7 a_1184_n1432# a_1184_1000# a_n2126_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_J2NVFM a_n406_1000# a_n406_n1432# a_124_n1432#
+ a_124_1000# a_n536_n1562#
X0 a_124_n1432# a_124_1000# a_n536_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X1 a_n406_n1432# a_n406_1000# a_n536_n1562# sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
.ends

.subckt isource_conv m1_4090_13100# m1_9600_7000# m1_4700_7820# m2_10060_7720# m1_5350_12620#
+ sky130_fd_pr__res_xhigh_po_1p41_BQY2W7_0/a_1714_n1432# li_9700_9140# VSUBS m1_4150_7820#
Xisource_cmirror_0 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_1 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_2 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_3 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_4 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xisource_cmirror_5 m1_9600_7000# li_9700_9140# m2_10060_7720# m1_5350_12620# isource_cmirror
Xsky130_fd_pr__res_xhigh_po_1p41_BQY2W7_0 m1_6360_10260# m1_5300_10260# m1_4700_7820#
+ m1_7960_7820# m1_8480_10260# sky130_fd_pr__res_xhigh_po_1p41_BQY2W7_0/a_1714_n1432#
+ m1_7960_7820# m1_5300_10260# m1_8480_10260# VSUBS m1_6900_7820# m1_7420_10260# m1_6360_10260#
+ m1_5840_7820# m1_5840_7820# m1_6900_7820# m1_7420_10260# sky130_fd_pr__res_xhigh_po_1p41_BQY2W7
Xsky130_fd_pr__nfet_01v8_WY4VMC_2 m1_5350_12620# m1_4090_13100# m1_4150_7820# VSUBS
+ m1_4090_13100# m1_4150_7820# sky130_fd_pr__nfet_01v8_WY4VMC
Xsky130_fd_pr__res_xhigh_po_1p41_J2NVFM_0 m1_4160_10260# m1_4150_7820# m1_4700_7820#
+ m1_4160_10260# VSUBS sky130_fd_pr__res_xhigh_po_1p41_J2NVFM
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ZZ3Y87 a_n287_n909# a_n229_n997# a_n1003_n997#
+ a_229_109# a_n1061_n909# a_287_n997# a_n487_21# a_n1061_109# a_745_n909# a_n545_109#
+ a_287_21# a_n1261_21# a_1061_n997# a_487_109# a_n745_21# a_229_n909# a_n29_109#
+ a_1061_21# a_29_21# a_n487_n997# a_n1261_n997# a_545_21# a_n545_n909# a_n287_109#
+ a_545_n997# a_1003_n909# a_1003_109# a_n29_n909# a_803_21# a_487_n909# a_29_n997#
+ a_n229_21# a_n745_n997# a_n803_n909# a_n803_109# a_n1319_109# a_803_n997# a_1261_109#
+ a_n1003_21# a_n1421_n1083# a_1261_n909# a_745_109# a_n1319_n909#
X0 a_229_109# a_29_21# a_n29_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X1 a_1261_n909# a_1061_n997# a_1003_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X2 a_487_109# a_287_21# a_229_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=1e+06u
X3 a_n545_109# a_n745_21# a_n803_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X4 a_1261_109# a_1061_21# a_1003_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X5 a_n29_n909# a_n229_n997# a_n287_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X6 a_229_n909# a_29_n997# a_n29_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=1e+06u
X7 a_n1061_109# a_n1261_21# a_n1319_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X8 a_n287_109# a_n487_21# a_n545_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=1e+06u
X9 a_n545_n909# a_n745_n997# a_n803_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X10 a_n287_n909# a_n487_n997# a_n545_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X11 a_n803_n909# a_n1003_n997# a_n1061_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X12 a_1003_109# a_803_21# a_745_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X13 a_n1061_n909# a_n1261_n997# a_n1319_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X14 a_1003_n909# a_803_n997# a_745_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X15 a_n803_109# a_n1003_21# a_n1061_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X16 a_745_n909# a_545_n997# a_487_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X17 a_n29_109# a_n229_21# a_n287_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X18 a_745_109# a_545_21# a_487_109# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X19 a_487_n909# a_287_n997# a_229_n909# a_n1421_n1083# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
.ends

.subckt isource_diffamp dw_14640_n8120# w_14846_n7914# m1_15050_n7600# m1_14640_n6760#
+ m1_15310_n7040#
Xsky130_fd_pr__nfet_01v8_lvt_ZZ3Y87_0 m1_15050_n7600# m1_14640_n6760# m1_14640_n6760#
+ m1_15050_n7600# m1_15310_n7040# m1_14640_n6760# m1_14640_n6760# m1_15310_n7040#
+ m1_15050_n7600# m1_15310_n7040# m1_14640_n6760# m1_14640_n6760# m1_14640_n6760#
+ m1_15310_n7040# m1_14640_n6760# m1_15050_n7600# m1_15310_n7040# m1_14640_n6760#
+ m1_14640_n6760# m1_14640_n6760# m1_14640_n6760# m1_14640_n6760# m1_15310_n7040#
+ m1_15050_n7600# m1_14640_n6760# m1_15310_n7040# m1_15310_n7040# m1_15310_n7040#
+ m1_14640_n6760# m1_15310_n7040# m1_14640_n6760# m1_14640_n6760# m1_14640_n6760#
+ m1_15050_n7600# m1_15050_n7600# m1_15050_n7600# m1_14640_n6760# m1_15050_n7600#
+ m1_14640_n6760# w_14846_n7914# m1_15050_n7600# m1_15050_n7600# m1_15050_n7600# sky130_fd_pr__nfet_01v8_lvt_ZZ3Y87
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG#1 m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt isource VP I_ref VM12G VM11D VN VM2D
Xsky130_fd_pr__cap_mim_m3_1_WXTTNJ_0 VP VM8D sky130_fd_pr__cap_mim_m3_1_WXTTNJ#0
Xisource_out_0 VM3D VM8D VM3G VM22D VP VN I_ref isource_out
Xisource_conv_tsmal_nwell_0 VP VM12G VM12G VP VM14D isource_conv_tsmal_nwell
Xisource_startup_0 VP VM11D VM8D VN isource_startup
Xisource_ref_0 VM11D VM11D VM12G VM2D VM12D VN isource_ref
Xisource_cmirror_2 VM8D VP VM9D isource_cmirror#0
Xisource_cmirror_3 VM8D VP VM8D isource_cmirror#0
Xisource_conv_0 VN VM8D VM3G m2_19160_1520# VM14D VN VP VN VM12G isource_conv
Xisource_diffamp_0 VP VM11D VM11D VM9D VM8D isource_diffamp
Xisource_diffamp_1 VP VM2D VM2D VM9D VM9D isource_diffamp
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_0 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#1
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_1 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#1
.ends


Xcurr_mirror_distribution_0 VP isource_0/I_ref curr_mirror_channel_0/I_in curr_mirror_distribution
Xtia_core_0 VP tia_core_0/Out_2 comparator_0/In tia_core_0/Disable_TIA tia_core_0/I_Bias1
+ outd_0/InputRef tia_core_0/VM39D tia_core_0/Input VN tia_core
Xtransmitter_0 VN curr_mirror_channel_0/LVDS_Bias transmitter_0/In transmitter
Xoutd_0 VP outd_0/InputRef outd_0/I_Bias outd_0/outd_stage1_0/isource_out outd_0/VM1_D
+ outd_0/VM14D comparator_0/In VN outd
Xcurr_mirror_channel_0 tia_core_0/I_Bias1 curr_mirror_channel_0/Comp_Bias_6 curr_mirror_channel_0/Comp_Bias_5
+ curr_mirror_channel_0/ctl_Bias VP curr_mirror_channel_0/Comp_Bias_3 curr_mirror_channel_0/Comp_Bias_2
+ curr_mirror_channel_0/Comp_Bias_1 curr_mirror_channel_0/LVDS_Bias curr_mirror_channel_0/I_in
+ comparator_0/comp_adv3_2/bias outd_0/I_Bias VN curr_mirror_channel
Xcomparator_0 curr_mirror_channel_0/Comp_Bias_6 VP comparator_0/comp_adv3_2/bias curr_mirror_channel_0/Comp_Bias_3
+ outd_0/InputRef curr_mirror_channel_0/ctl_Bias curr_mirror_channel_0/Comp_Bias_5
+ transmitter_0/In comparator_0/In VN comparator
Xfb_dark_current_0 VP comparator_0/In outd_0/InputRef VN fb_dark_current
Xisource_0 VP isource_0/I_ref isource_0/VM12G isource_0/VM11D VN isource_0/VM2D isource


