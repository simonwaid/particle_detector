magic
tech sky130B
magscale 1 2
timestamp 1654605132
<< error_p >>
rect -365 1508 -307 1514
rect -173 1508 -115 1514
rect 19 1508 77 1514
rect 211 1508 269 1514
rect 403 1508 461 1514
rect -365 1474 -353 1508
rect -173 1474 -161 1508
rect 19 1474 31 1508
rect 211 1474 223 1508
rect 403 1474 415 1508
rect -365 1468 -307 1474
rect -173 1468 -115 1474
rect 19 1468 77 1474
rect 211 1468 269 1474
rect 403 1468 461 1474
rect -461 998 -403 1004
rect -269 998 -211 1004
rect -77 998 -19 1004
rect 115 998 173 1004
rect 307 998 365 1004
rect -461 964 -449 998
rect -269 964 -257 998
rect -77 964 -65 998
rect 115 964 127 998
rect 307 964 319 998
rect -461 958 -403 964
rect -269 958 -211 964
rect -77 958 -19 964
rect 115 958 173 964
rect 307 958 365 964
rect -461 890 -403 896
rect -269 890 -211 896
rect -77 890 -19 896
rect 115 890 173 896
rect 307 890 365 896
rect -461 856 -449 890
rect -269 856 -257 890
rect -77 856 -65 890
rect 115 856 127 890
rect 307 856 319 890
rect -461 850 -403 856
rect -269 850 -211 856
rect -77 850 -19 856
rect 115 850 173 856
rect 307 850 365 856
rect -365 380 -307 386
rect -173 380 -115 386
rect 19 380 77 386
rect 211 380 269 386
rect 403 380 461 386
rect -365 346 -353 380
rect -173 346 -161 380
rect 19 346 31 380
rect 211 346 223 380
rect 403 346 415 380
rect -365 340 -307 346
rect -173 340 -115 346
rect 19 340 77 346
rect 211 340 269 346
rect 403 340 461 346
rect -365 272 -307 278
rect -173 272 -115 278
rect 19 272 77 278
rect 211 272 269 278
rect 403 272 461 278
rect -365 238 -353 272
rect -173 238 -161 272
rect 19 238 31 272
rect 211 238 223 272
rect 403 238 415 272
rect -365 232 -307 238
rect -173 232 -115 238
rect 19 232 77 238
rect 211 232 269 238
rect 403 232 461 238
rect -461 -238 -403 -232
rect -269 -238 -211 -232
rect -77 -238 -19 -232
rect 115 -238 173 -232
rect 307 -238 365 -232
rect -461 -272 -449 -238
rect -269 -272 -257 -238
rect -77 -272 -65 -238
rect 115 -272 127 -238
rect 307 -272 319 -238
rect -461 -278 -403 -272
rect -269 -278 -211 -272
rect -77 -278 -19 -272
rect 115 -278 173 -272
rect 307 -278 365 -272
rect -461 -346 -403 -340
rect -269 -346 -211 -340
rect -77 -346 -19 -340
rect 115 -346 173 -340
rect 307 -346 365 -340
rect -461 -380 -449 -346
rect -269 -380 -257 -346
rect -77 -380 -65 -346
rect 115 -380 127 -346
rect 307 -380 319 -346
rect -461 -386 -403 -380
rect -269 -386 -211 -380
rect -77 -386 -19 -380
rect 115 -386 173 -380
rect 307 -386 365 -380
rect -365 -856 -307 -850
rect -173 -856 -115 -850
rect 19 -856 77 -850
rect 211 -856 269 -850
rect 403 -856 461 -850
rect -365 -890 -353 -856
rect -173 -890 -161 -856
rect 19 -890 31 -856
rect 211 -890 223 -856
rect 403 -890 415 -856
rect -365 -896 -307 -890
rect -173 -896 -115 -890
rect 19 -896 77 -890
rect 211 -896 269 -890
rect 403 -896 461 -890
rect -365 -964 -307 -958
rect -173 -964 -115 -958
rect 19 -964 77 -958
rect 211 -964 269 -958
rect 403 -964 461 -958
rect -365 -998 -353 -964
rect -173 -998 -161 -964
rect 19 -998 31 -964
rect 211 -998 223 -964
rect 403 -998 415 -964
rect -365 -1004 -307 -998
rect -173 -1004 -115 -998
rect 19 -1004 77 -998
rect 211 -1004 269 -998
rect 403 -1004 461 -998
rect -461 -1474 -403 -1468
rect -269 -1474 -211 -1468
rect -77 -1474 -19 -1468
rect 115 -1474 173 -1468
rect 307 -1474 365 -1468
rect -461 -1508 -449 -1474
rect -269 -1508 -257 -1474
rect -77 -1508 -65 -1474
rect 115 -1508 127 -1474
rect 307 -1508 319 -1474
rect -461 -1514 -403 -1508
rect -269 -1514 -211 -1508
rect -77 -1514 -19 -1508
rect 115 -1514 173 -1508
rect 307 -1514 365 -1508
<< pwell >>
rect -647 -1646 647 1646
<< nmoslvt >>
rect -447 1036 -417 1436
rect -351 1036 -321 1436
rect -255 1036 -225 1436
rect -159 1036 -129 1436
rect -63 1036 -33 1436
rect 33 1036 63 1436
rect 129 1036 159 1436
rect 225 1036 255 1436
rect 321 1036 351 1436
rect 417 1036 447 1436
rect -447 418 -417 818
rect -351 418 -321 818
rect -255 418 -225 818
rect -159 418 -129 818
rect -63 418 -33 818
rect 33 418 63 818
rect 129 418 159 818
rect 225 418 255 818
rect 321 418 351 818
rect 417 418 447 818
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect -447 -818 -417 -418
rect -351 -818 -321 -418
rect -255 -818 -225 -418
rect -159 -818 -129 -418
rect -63 -818 -33 -418
rect 33 -818 63 -418
rect 129 -818 159 -418
rect 225 -818 255 -418
rect 321 -818 351 -418
rect 417 -818 447 -418
rect -447 -1436 -417 -1036
rect -351 -1436 -321 -1036
rect -255 -1436 -225 -1036
rect -159 -1436 -129 -1036
rect -63 -1436 -33 -1036
rect 33 -1436 63 -1036
rect 129 -1436 159 -1036
rect 225 -1436 255 -1036
rect 321 -1436 351 -1036
rect 417 -1436 447 -1036
<< ndiff >>
rect -509 1424 -447 1436
rect -509 1048 -497 1424
rect -463 1048 -447 1424
rect -509 1036 -447 1048
rect -417 1424 -351 1436
rect -417 1048 -401 1424
rect -367 1048 -351 1424
rect -417 1036 -351 1048
rect -321 1424 -255 1436
rect -321 1048 -305 1424
rect -271 1048 -255 1424
rect -321 1036 -255 1048
rect -225 1424 -159 1436
rect -225 1048 -209 1424
rect -175 1048 -159 1424
rect -225 1036 -159 1048
rect -129 1424 -63 1436
rect -129 1048 -113 1424
rect -79 1048 -63 1424
rect -129 1036 -63 1048
rect -33 1424 33 1436
rect -33 1048 -17 1424
rect 17 1048 33 1424
rect -33 1036 33 1048
rect 63 1424 129 1436
rect 63 1048 79 1424
rect 113 1048 129 1424
rect 63 1036 129 1048
rect 159 1424 225 1436
rect 159 1048 175 1424
rect 209 1048 225 1424
rect 159 1036 225 1048
rect 255 1424 321 1436
rect 255 1048 271 1424
rect 305 1048 321 1424
rect 255 1036 321 1048
rect 351 1424 417 1436
rect 351 1048 367 1424
rect 401 1048 417 1424
rect 351 1036 417 1048
rect 447 1424 509 1436
rect 447 1048 463 1424
rect 497 1048 509 1424
rect 447 1036 509 1048
rect -509 806 -447 818
rect -509 430 -497 806
rect -463 430 -447 806
rect -509 418 -447 430
rect -417 806 -351 818
rect -417 430 -401 806
rect -367 430 -351 806
rect -417 418 -351 430
rect -321 806 -255 818
rect -321 430 -305 806
rect -271 430 -255 806
rect -321 418 -255 430
rect -225 806 -159 818
rect -225 430 -209 806
rect -175 430 -159 806
rect -225 418 -159 430
rect -129 806 -63 818
rect -129 430 -113 806
rect -79 430 -63 806
rect -129 418 -63 430
rect -33 806 33 818
rect -33 430 -17 806
rect 17 430 33 806
rect -33 418 33 430
rect 63 806 129 818
rect 63 430 79 806
rect 113 430 129 806
rect 63 418 129 430
rect 159 806 225 818
rect 159 430 175 806
rect 209 430 225 806
rect 159 418 225 430
rect 255 806 321 818
rect 255 430 271 806
rect 305 430 321 806
rect 255 418 321 430
rect 351 806 417 818
rect 351 430 367 806
rect 401 430 417 806
rect 351 418 417 430
rect 447 806 509 818
rect 447 430 463 806
rect 497 430 509 806
rect 447 418 509 430
rect -509 188 -447 200
rect -509 -188 -497 188
rect -463 -188 -447 188
rect -509 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 509 200
rect 447 -188 463 188
rect 497 -188 509 188
rect 447 -200 509 -188
rect -509 -430 -447 -418
rect -509 -806 -497 -430
rect -463 -806 -447 -430
rect -509 -818 -447 -806
rect -417 -430 -351 -418
rect -417 -806 -401 -430
rect -367 -806 -351 -430
rect -417 -818 -351 -806
rect -321 -430 -255 -418
rect -321 -806 -305 -430
rect -271 -806 -255 -430
rect -321 -818 -255 -806
rect -225 -430 -159 -418
rect -225 -806 -209 -430
rect -175 -806 -159 -430
rect -225 -818 -159 -806
rect -129 -430 -63 -418
rect -129 -806 -113 -430
rect -79 -806 -63 -430
rect -129 -818 -63 -806
rect -33 -430 33 -418
rect -33 -806 -17 -430
rect 17 -806 33 -430
rect -33 -818 33 -806
rect 63 -430 129 -418
rect 63 -806 79 -430
rect 113 -806 129 -430
rect 63 -818 129 -806
rect 159 -430 225 -418
rect 159 -806 175 -430
rect 209 -806 225 -430
rect 159 -818 225 -806
rect 255 -430 321 -418
rect 255 -806 271 -430
rect 305 -806 321 -430
rect 255 -818 321 -806
rect 351 -430 417 -418
rect 351 -806 367 -430
rect 401 -806 417 -430
rect 351 -818 417 -806
rect 447 -430 509 -418
rect 447 -806 463 -430
rect 497 -806 509 -430
rect 447 -818 509 -806
rect -509 -1048 -447 -1036
rect -509 -1424 -497 -1048
rect -463 -1424 -447 -1048
rect -509 -1436 -447 -1424
rect -417 -1048 -351 -1036
rect -417 -1424 -401 -1048
rect -367 -1424 -351 -1048
rect -417 -1436 -351 -1424
rect -321 -1048 -255 -1036
rect -321 -1424 -305 -1048
rect -271 -1424 -255 -1048
rect -321 -1436 -255 -1424
rect -225 -1048 -159 -1036
rect -225 -1424 -209 -1048
rect -175 -1424 -159 -1048
rect -225 -1436 -159 -1424
rect -129 -1048 -63 -1036
rect -129 -1424 -113 -1048
rect -79 -1424 -63 -1048
rect -129 -1436 -63 -1424
rect -33 -1048 33 -1036
rect -33 -1424 -17 -1048
rect 17 -1424 33 -1048
rect -33 -1436 33 -1424
rect 63 -1048 129 -1036
rect 63 -1424 79 -1048
rect 113 -1424 129 -1048
rect 63 -1436 129 -1424
rect 159 -1048 225 -1036
rect 159 -1424 175 -1048
rect 209 -1424 225 -1048
rect 159 -1436 225 -1424
rect 255 -1048 321 -1036
rect 255 -1424 271 -1048
rect 305 -1424 321 -1048
rect 255 -1436 321 -1424
rect 351 -1048 417 -1036
rect 351 -1424 367 -1048
rect 401 -1424 417 -1048
rect 351 -1436 417 -1424
rect 447 -1048 509 -1036
rect 447 -1424 463 -1048
rect 497 -1424 509 -1048
rect 447 -1436 509 -1424
<< ndiffc >>
rect -497 1048 -463 1424
rect -401 1048 -367 1424
rect -305 1048 -271 1424
rect -209 1048 -175 1424
rect -113 1048 -79 1424
rect -17 1048 17 1424
rect 79 1048 113 1424
rect 175 1048 209 1424
rect 271 1048 305 1424
rect 367 1048 401 1424
rect 463 1048 497 1424
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect -497 -1424 -463 -1048
rect -401 -1424 -367 -1048
rect -305 -1424 -271 -1048
rect -209 -1424 -175 -1048
rect -113 -1424 -79 -1048
rect -17 -1424 17 -1048
rect 79 -1424 113 -1048
rect 175 -1424 209 -1048
rect 271 -1424 305 -1048
rect 367 -1424 401 -1048
rect 463 -1424 497 -1048
<< psubdiff >>
rect -611 1576 -515 1610
rect 515 1576 611 1610
rect -611 1514 -577 1576
rect 577 1514 611 1576
rect -611 -1576 -577 -1514
rect 577 -1576 611 -1514
rect -611 -1610 -515 -1576
rect 515 -1610 611 -1576
<< psubdiffcont >>
rect -515 1576 515 1610
rect -611 -1514 -577 1514
rect 577 -1514 611 1514
rect -515 -1610 515 -1576
<< poly >>
rect -369 1508 -303 1524
rect -369 1474 -353 1508
rect -319 1474 -303 1508
rect -447 1436 -417 1462
rect -369 1458 -303 1474
rect -177 1508 -111 1524
rect -177 1474 -161 1508
rect -127 1474 -111 1508
rect -351 1436 -321 1458
rect -255 1436 -225 1462
rect -177 1458 -111 1474
rect 15 1508 81 1524
rect 15 1474 31 1508
rect 65 1474 81 1508
rect -159 1436 -129 1458
rect -63 1436 -33 1462
rect 15 1458 81 1474
rect 207 1508 273 1524
rect 207 1474 223 1508
rect 257 1474 273 1508
rect 33 1436 63 1458
rect 129 1436 159 1462
rect 207 1458 273 1474
rect 399 1508 465 1524
rect 399 1474 415 1508
rect 449 1474 465 1508
rect 225 1436 255 1458
rect 321 1436 351 1462
rect 399 1458 465 1474
rect 417 1436 447 1458
rect -447 1014 -417 1036
rect -465 998 -399 1014
rect -351 1010 -321 1036
rect -255 1014 -225 1036
rect -465 964 -449 998
rect -415 964 -399 998
rect -465 948 -399 964
rect -273 998 -207 1014
rect -159 1010 -129 1036
rect -63 1014 -33 1036
rect -273 964 -257 998
rect -223 964 -207 998
rect -273 948 -207 964
rect -81 998 -15 1014
rect 33 1010 63 1036
rect 129 1014 159 1036
rect -81 964 -65 998
rect -31 964 -15 998
rect -81 948 -15 964
rect 111 998 177 1014
rect 225 1010 255 1036
rect 321 1014 351 1036
rect 111 964 127 998
rect 161 964 177 998
rect 111 948 177 964
rect 303 998 369 1014
rect 417 1010 447 1036
rect 303 964 319 998
rect 353 964 369 998
rect 303 948 369 964
rect -465 890 -399 906
rect -465 856 -449 890
rect -415 856 -399 890
rect -465 840 -399 856
rect -273 890 -207 906
rect -273 856 -257 890
rect -223 856 -207 890
rect -447 818 -417 840
rect -351 818 -321 844
rect -273 840 -207 856
rect -81 890 -15 906
rect -81 856 -65 890
rect -31 856 -15 890
rect -255 818 -225 840
rect -159 818 -129 844
rect -81 840 -15 856
rect 111 890 177 906
rect 111 856 127 890
rect 161 856 177 890
rect -63 818 -33 840
rect 33 818 63 844
rect 111 840 177 856
rect 303 890 369 906
rect 303 856 319 890
rect 353 856 369 890
rect 129 818 159 840
rect 225 818 255 844
rect 303 840 369 856
rect 321 818 351 840
rect 417 818 447 844
rect -447 392 -417 418
rect -351 396 -321 418
rect -369 380 -303 396
rect -255 392 -225 418
rect -159 396 -129 418
rect -369 346 -353 380
rect -319 346 -303 380
rect -369 330 -303 346
rect -177 380 -111 396
rect -63 392 -33 418
rect 33 396 63 418
rect -177 346 -161 380
rect -127 346 -111 380
rect -177 330 -111 346
rect 15 380 81 396
rect 129 392 159 418
rect 225 396 255 418
rect 15 346 31 380
rect 65 346 81 380
rect 15 330 81 346
rect 207 380 273 396
rect 321 392 351 418
rect 417 396 447 418
rect 207 346 223 380
rect 257 346 273 380
rect 207 330 273 346
rect 399 380 465 396
rect 399 346 415 380
rect 449 346 465 380
rect 399 330 465 346
rect -369 272 -303 288
rect -369 238 -353 272
rect -319 238 -303 272
rect -447 200 -417 226
rect -369 222 -303 238
rect -177 272 -111 288
rect -177 238 -161 272
rect -127 238 -111 272
rect -351 200 -321 222
rect -255 200 -225 226
rect -177 222 -111 238
rect 15 272 81 288
rect 15 238 31 272
rect 65 238 81 272
rect -159 200 -129 222
rect -63 200 -33 226
rect 15 222 81 238
rect 207 272 273 288
rect 207 238 223 272
rect 257 238 273 272
rect 33 200 63 222
rect 129 200 159 226
rect 207 222 273 238
rect 399 272 465 288
rect 399 238 415 272
rect 449 238 465 272
rect 225 200 255 222
rect 321 200 351 226
rect 399 222 465 238
rect 417 200 447 222
rect -447 -222 -417 -200
rect -465 -238 -399 -222
rect -351 -226 -321 -200
rect -255 -222 -225 -200
rect -465 -272 -449 -238
rect -415 -272 -399 -238
rect -465 -288 -399 -272
rect -273 -238 -207 -222
rect -159 -226 -129 -200
rect -63 -222 -33 -200
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -273 -288 -207 -272
rect -81 -238 -15 -222
rect 33 -226 63 -200
rect 129 -222 159 -200
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect -81 -288 -15 -272
rect 111 -238 177 -222
rect 225 -226 255 -200
rect 321 -222 351 -200
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 111 -288 177 -272
rect 303 -238 369 -222
rect 417 -226 447 -200
rect 303 -272 319 -238
rect 353 -272 369 -238
rect 303 -288 369 -272
rect -465 -346 -399 -330
rect -465 -380 -449 -346
rect -415 -380 -399 -346
rect -465 -396 -399 -380
rect -273 -346 -207 -330
rect -273 -380 -257 -346
rect -223 -380 -207 -346
rect -447 -418 -417 -396
rect -351 -418 -321 -392
rect -273 -396 -207 -380
rect -81 -346 -15 -330
rect -81 -380 -65 -346
rect -31 -380 -15 -346
rect -255 -418 -225 -396
rect -159 -418 -129 -392
rect -81 -396 -15 -380
rect 111 -346 177 -330
rect 111 -380 127 -346
rect 161 -380 177 -346
rect -63 -418 -33 -396
rect 33 -418 63 -392
rect 111 -396 177 -380
rect 303 -346 369 -330
rect 303 -380 319 -346
rect 353 -380 369 -346
rect 129 -418 159 -396
rect 225 -418 255 -392
rect 303 -396 369 -380
rect 321 -418 351 -396
rect 417 -418 447 -392
rect -447 -844 -417 -818
rect -351 -840 -321 -818
rect -369 -856 -303 -840
rect -255 -844 -225 -818
rect -159 -840 -129 -818
rect -369 -890 -353 -856
rect -319 -890 -303 -856
rect -369 -906 -303 -890
rect -177 -856 -111 -840
rect -63 -844 -33 -818
rect 33 -840 63 -818
rect -177 -890 -161 -856
rect -127 -890 -111 -856
rect -177 -906 -111 -890
rect 15 -856 81 -840
rect 129 -844 159 -818
rect 225 -840 255 -818
rect 15 -890 31 -856
rect 65 -890 81 -856
rect 15 -906 81 -890
rect 207 -856 273 -840
rect 321 -844 351 -818
rect 417 -840 447 -818
rect 207 -890 223 -856
rect 257 -890 273 -856
rect 207 -906 273 -890
rect 399 -856 465 -840
rect 399 -890 415 -856
rect 449 -890 465 -856
rect 399 -906 465 -890
rect -369 -964 -303 -948
rect -369 -998 -353 -964
rect -319 -998 -303 -964
rect -447 -1036 -417 -1010
rect -369 -1014 -303 -998
rect -177 -964 -111 -948
rect -177 -998 -161 -964
rect -127 -998 -111 -964
rect -351 -1036 -321 -1014
rect -255 -1036 -225 -1010
rect -177 -1014 -111 -998
rect 15 -964 81 -948
rect 15 -998 31 -964
rect 65 -998 81 -964
rect -159 -1036 -129 -1014
rect -63 -1036 -33 -1010
rect 15 -1014 81 -998
rect 207 -964 273 -948
rect 207 -998 223 -964
rect 257 -998 273 -964
rect 33 -1036 63 -1014
rect 129 -1036 159 -1010
rect 207 -1014 273 -998
rect 399 -964 465 -948
rect 399 -998 415 -964
rect 449 -998 465 -964
rect 225 -1036 255 -1014
rect 321 -1036 351 -1010
rect 399 -1014 465 -998
rect 417 -1036 447 -1014
rect -447 -1458 -417 -1436
rect -465 -1474 -399 -1458
rect -351 -1462 -321 -1436
rect -255 -1458 -225 -1436
rect -465 -1508 -449 -1474
rect -415 -1508 -399 -1474
rect -465 -1524 -399 -1508
rect -273 -1474 -207 -1458
rect -159 -1462 -129 -1436
rect -63 -1458 -33 -1436
rect -273 -1508 -257 -1474
rect -223 -1508 -207 -1474
rect -273 -1524 -207 -1508
rect -81 -1474 -15 -1458
rect 33 -1462 63 -1436
rect 129 -1458 159 -1436
rect -81 -1508 -65 -1474
rect -31 -1508 -15 -1474
rect -81 -1524 -15 -1508
rect 111 -1474 177 -1458
rect 225 -1462 255 -1436
rect 321 -1458 351 -1436
rect 111 -1508 127 -1474
rect 161 -1508 177 -1474
rect 111 -1524 177 -1508
rect 303 -1474 369 -1458
rect 417 -1462 447 -1436
rect 303 -1508 319 -1474
rect 353 -1508 369 -1474
rect 303 -1524 369 -1508
<< polycont >>
rect -353 1474 -319 1508
rect -161 1474 -127 1508
rect 31 1474 65 1508
rect 223 1474 257 1508
rect 415 1474 449 1508
rect -449 964 -415 998
rect -257 964 -223 998
rect -65 964 -31 998
rect 127 964 161 998
rect 319 964 353 998
rect -449 856 -415 890
rect -257 856 -223 890
rect -65 856 -31 890
rect 127 856 161 890
rect 319 856 353 890
rect -353 346 -319 380
rect -161 346 -127 380
rect 31 346 65 380
rect 223 346 257 380
rect 415 346 449 380
rect -353 238 -319 272
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect 415 238 449 272
rect -449 -272 -415 -238
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
rect 319 -272 353 -238
rect -449 -380 -415 -346
rect -257 -380 -223 -346
rect -65 -380 -31 -346
rect 127 -380 161 -346
rect 319 -380 353 -346
rect -353 -890 -319 -856
rect -161 -890 -127 -856
rect 31 -890 65 -856
rect 223 -890 257 -856
rect 415 -890 449 -856
rect -353 -998 -319 -964
rect -161 -998 -127 -964
rect 31 -998 65 -964
rect 223 -998 257 -964
rect 415 -998 449 -964
rect -449 -1508 -415 -1474
rect -257 -1508 -223 -1474
rect -65 -1508 -31 -1474
rect 127 -1508 161 -1474
rect 319 -1508 353 -1474
<< locali >>
rect -611 1576 -515 1610
rect 515 1576 611 1610
rect -611 1514 -577 1576
rect 577 1514 611 1576
rect -369 1474 -353 1508
rect -319 1474 -303 1508
rect -177 1474 -161 1508
rect -127 1474 -111 1508
rect 15 1474 31 1508
rect 65 1474 81 1508
rect 207 1474 223 1508
rect 257 1474 273 1508
rect 399 1474 415 1508
rect 449 1474 465 1508
rect -497 1424 -463 1440
rect -497 1032 -463 1048
rect -401 1424 -367 1440
rect -401 1032 -367 1048
rect -305 1424 -271 1440
rect -305 1032 -271 1048
rect -209 1424 -175 1440
rect -209 1032 -175 1048
rect -113 1424 -79 1440
rect -113 1032 -79 1048
rect -17 1424 17 1440
rect -17 1032 17 1048
rect 79 1424 113 1440
rect 79 1032 113 1048
rect 175 1424 209 1440
rect 175 1032 209 1048
rect 271 1424 305 1440
rect 271 1032 305 1048
rect 367 1424 401 1440
rect 367 1032 401 1048
rect 463 1424 497 1440
rect 463 1032 497 1048
rect -465 964 -449 998
rect -415 964 -399 998
rect -273 964 -257 998
rect -223 964 -207 998
rect -81 964 -65 998
rect -31 964 -15 998
rect 111 964 127 998
rect 161 964 177 998
rect 303 964 319 998
rect 353 964 369 998
rect -465 856 -449 890
rect -415 856 -399 890
rect -273 856 -257 890
rect -223 856 -207 890
rect -81 856 -65 890
rect -31 856 -15 890
rect 111 856 127 890
rect 161 856 177 890
rect 303 856 319 890
rect 353 856 369 890
rect -497 806 -463 822
rect -497 414 -463 430
rect -401 806 -367 822
rect -401 414 -367 430
rect -305 806 -271 822
rect -305 414 -271 430
rect -209 806 -175 822
rect -209 414 -175 430
rect -113 806 -79 822
rect -113 414 -79 430
rect -17 806 17 822
rect -17 414 17 430
rect 79 806 113 822
rect 79 414 113 430
rect 175 806 209 822
rect 175 414 209 430
rect 271 806 305 822
rect 271 414 305 430
rect 367 806 401 822
rect 367 414 401 430
rect 463 806 497 822
rect 463 414 497 430
rect -369 346 -353 380
rect -319 346 -303 380
rect -177 346 -161 380
rect -127 346 -111 380
rect 15 346 31 380
rect 65 346 81 380
rect 207 346 223 380
rect 257 346 273 380
rect 399 346 415 380
rect 449 346 465 380
rect -369 238 -353 272
rect -319 238 -303 272
rect -177 238 -161 272
rect -127 238 -111 272
rect 15 238 31 272
rect 65 238 81 272
rect 207 238 223 272
rect 257 238 273 272
rect 399 238 415 272
rect 449 238 465 272
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect -465 -272 -449 -238
rect -415 -272 -399 -238
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 303 -272 319 -238
rect 353 -272 369 -238
rect -465 -380 -449 -346
rect -415 -380 -399 -346
rect -273 -380 -257 -346
rect -223 -380 -207 -346
rect -81 -380 -65 -346
rect -31 -380 -15 -346
rect 111 -380 127 -346
rect 161 -380 177 -346
rect 303 -380 319 -346
rect 353 -380 369 -346
rect -497 -430 -463 -414
rect -497 -822 -463 -806
rect -401 -430 -367 -414
rect -401 -822 -367 -806
rect -305 -430 -271 -414
rect -305 -822 -271 -806
rect -209 -430 -175 -414
rect -209 -822 -175 -806
rect -113 -430 -79 -414
rect -113 -822 -79 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 79 -430 113 -414
rect 79 -822 113 -806
rect 175 -430 209 -414
rect 175 -822 209 -806
rect 271 -430 305 -414
rect 271 -822 305 -806
rect 367 -430 401 -414
rect 367 -822 401 -806
rect 463 -430 497 -414
rect 463 -822 497 -806
rect -369 -890 -353 -856
rect -319 -890 -303 -856
rect -177 -890 -161 -856
rect -127 -890 -111 -856
rect 15 -890 31 -856
rect 65 -890 81 -856
rect 207 -890 223 -856
rect 257 -890 273 -856
rect 399 -890 415 -856
rect 449 -890 465 -856
rect -369 -998 -353 -964
rect -319 -998 -303 -964
rect -177 -998 -161 -964
rect -127 -998 -111 -964
rect 15 -998 31 -964
rect 65 -998 81 -964
rect 207 -998 223 -964
rect 257 -998 273 -964
rect 399 -998 415 -964
rect 449 -998 465 -964
rect -497 -1048 -463 -1032
rect -497 -1440 -463 -1424
rect -401 -1048 -367 -1032
rect -401 -1440 -367 -1424
rect -305 -1048 -271 -1032
rect -305 -1440 -271 -1424
rect -209 -1048 -175 -1032
rect -209 -1440 -175 -1424
rect -113 -1048 -79 -1032
rect -113 -1440 -79 -1424
rect -17 -1048 17 -1032
rect -17 -1440 17 -1424
rect 79 -1048 113 -1032
rect 79 -1440 113 -1424
rect 175 -1048 209 -1032
rect 175 -1440 209 -1424
rect 271 -1048 305 -1032
rect 271 -1440 305 -1424
rect 367 -1048 401 -1032
rect 367 -1440 401 -1424
rect 463 -1048 497 -1032
rect 463 -1440 497 -1424
rect -465 -1508 -449 -1474
rect -415 -1508 -399 -1474
rect -273 -1508 -257 -1474
rect -223 -1508 -207 -1474
rect -81 -1508 -65 -1474
rect -31 -1508 -15 -1474
rect 111 -1508 127 -1474
rect 161 -1508 177 -1474
rect 303 -1508 319 -1474
rect 353 -1508 369 -1474
rect -611 -1576 -577 -1514
rect 577 -1576 611 -1514
rect -611 -1610 -515 -1576
rect 515 -1610 611 -1576
<< viali >>
rect -353 1474 -319 1508
rect -161 1474 -127 1508
rect 31 1474 65 1508
rect 223 1474 257 1508
rect 415 1474 449 1508
rect -497 1048 -463 1424
rect -401 1048 -367 1424
rect -305 1048 -271 1424
rect -209 1048 -175 1424
rect -113 1048 -79 1424
rect -17 1048 17 1424
rect 79 1048 113 1424
rect 175 1048 209 1424
rect 271 1048 305 1424
rect 367 1048 401 1424
rect 463 1048 497 1424
rect -449 964 -415 998
rect -257 964 -223 998
rect -65 964 -31 998
rect 127 964 161 998
rect 319 964 353 998
rect -449 856 -415 890
rect -257 856 -223 890
rect -65 856 -31 890
rect 127 856 161 890
rect 319 856 353 890
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect -353 346 -319 380
rect -161 346 -127 380
rect 31 346 65 380
rect 223 346 257 380
rect 415 346 449 380
rect -353 238 -319 272
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect 415 238 449 272
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect -449 -272 -415 -238
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
rect 319 -272 353 -238
rect -449 -380 -415 -346
rect -257 -380 -223 -346
rect -65 -380 -31 -346
rect 127 -380 161 -346
rect 319 -380 353 -346
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect -353 -890 -319 -856
rect -161 -890 -127 -856
rect 31 -890 65 -856
rect 223 -890 257 -856
rect 415 -890 449 -856
rect -353 -998 -319 -964
rect -161 -998 -127 -964
rect 31 -998 65 -964
rect 223 -998 257 -964
rect 415 -998 449 -964
rect -497 -1424 -463 -1048
rect -401 -1424 -367 -1048
rect -305 -1424 -271 -1048
rect -209 -1424 -175 -1048
rect -113 -1424 -79 -1048
rect -17 -1424 17 -1048
rect 79 -1424 113 -1048
rect 175 -1424 209 -1048
rect 271 -1424 305 -1048
rect 367 -1424 401 -1048
rect 463 -1424 497 -1048
rect -449 -1508 -415 -1474
rect -257 -1508 -223 -1474
rect -65 -1508 -31 -1474
rect 127 -1508 161 -1474
rect 319 -1508 353 -1474
<< metal1 >>
rect -365 1508 -307 1514
rect -365 1474 -353 1508
rect -319 1474 -307 1508
rect -365 1468 -307 1474
rect -173 1508 -115 1514
rect -173 1474 -161 1508
rect -127 1474 -115 1508
rect -173 1468 -115 1474
rect 19 1508 77 1514
rect 19 1474 31 1508
rect 65 1474 77 1508
rect 19 1468 77 1474
rect 211 1508 269 1514
rect 211 1474 223 1508
rect 257 1474 269 1508
rect 211 1468 269 1474
rect 403 1508 461 1514
rect 403 1474 415 1508
rect 449 1474 461 1508
rect 403 1468 461 1474
rect -503 1424 -457 1436
rect -503 1048 -497 1424
rect -463 1048 -457 1424
rect -503 1036 -457 1048
rect -407 1424 -361 1436
rect -407 1048 -401 1424
rect -367 1048 -361 1424
rect -407 1036 -361 1048
rect -311 1424 -265 1436
rect -311 1048 -305 1424
rect -271 1048 -265 1424
rect -311 1036 -265 1048
rect -215 1424 -169 1436
rect -215 1048 -209 1424
rect -175 1048 -169 1424
rect -215 1036 -169 1048
rect -119 1424 -73 1436
rect -119 1048 -113 1424
rect -79 1048 -73 1424
rect -119 1036 -73 1048
rect -23 1424 23 1436
rect -23 1048 -17 1424
rect 17 1048 23 1424
rect -23 1036 23 1048
rect 73 1424 119 1436
rect 73 1048 79 1424
rect 113 1048 119 1424
rect 73 1036 119 1048
rect 169 1424 215 1436
rect 169 1048 175 1424
rect 209 1048 215 1424
rect 169 1036 215 1048
rect 265 1424 311 1436
rect 265 1048 271 1424
rect 305 1048 311 1424
rect 265 1036 311 1048
rect 361 1424 407 1436
rect 361 1048 367 1424
rect 401 1048 407 1424
rect 361 1036 407 1048
rect 457 1424 503 1436
rect 457 1048 463 1424
rect 497 1048 503 1424
rect 457 1036 503 1048
rect -461 998 -403 1004
rect -461 964 -449 998
rect -415 964 -403 998
rect -461 958 -403 964
rect -269 998 -211 1004
rect -269 964 -257 998
rect -223 964 -211 998
rect -269 958 -211 964
rect -77 998 -19 1004
rect -77 964 -65 998
rect -31 964 -19 998
rect -77 958 -19 964
rect 115 998 173 1004
rect 115 964 127 998
rect 161 964 173 998
rect 115 958 173 964
rect 307 998 365 1004
rect 307 964 319 998
rect 353 964 365 998
rect 307 958 365 964
rect -461 890 -403 896
rect -461 856 -449 890
rect -415 856 -403 890
rect -461 850 -403 856
rect -269 890 -211 896
rect -269 856 -257 890
rect -223 856 -211 890
rect -269 850 -211 856
rect -77 890 -19 896
rect -77 856 -65 890
rect -31 856 -19 890
rect -77 850 -19 856
rect 115 890 173 896
rect 115 856 127 890
rect 161 856 173 890
rect 115 850 173 856
rect 307 890 365 896
rect 307 856 319 890
rect 353 856 365 890
rect 307 850 365 856
rect -503 806 -457 818
rect -503 430 -497 806
rect -463 430 -457 806
rect -503 418 -457 430
rect -407 806 -361 818
rect -407 430 -401 806
rect -367 430 -361 806
rect -407 418 -361 430
rect -311 806 -265 818
rect -311 430 -305 806
rect -271 430 -265 806
rect -311 418 -265 430
rect -215 806 -169 818
rect -215 430 -209 806
rect -175 430 -169 806
rect -215 418 -169 430
rect -119 806 -73 818
rect -119 430 -113 806
rect -79 430 -73 806
rect -119 418 -73 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 73 806 119 818
rect 73 430 79 806
rect 113 430 119 806
rect 73 418 119 430
rect 169 806 215 818
rect 169 430 175 806
rect 209 430 215 806
rect 169 418 215 430
rect 265 806 311 818
rect 265 430 271 806
rect 305 430 311 806
rect 265 418 311 430
rect 361 806 407 818
rect 361 430 367 806
rect 401 430 407 806
rect 361 418 407 430
rect 457 806 503 818
rect 457 430 463 806
rect 497 430 503 806
rect 457 418 503 430
rect -365 380 -307 386
rect -365 346 -353 380
rect -319 346 -307 380
rect -365 340 -307 346
rect -173 380 -115 386
rect -173 346 -161 380
rect -127 346 -115 380
rect -173 340 -115 346
rect 19 380 77 386
rect 19 346 31 380
rect 65 346 77 380
rect 19 340 77 346
rect 211 380 269 386
rect 211 346 223 380
rect 257 346 269 380
rect 211 340 269 346
rect 403 380 461 386
rect 403 346 415 380
rect 449 346 461 380
rect 403 340 461 346
rect -365 272 -307 278
rect -365 238 -353 272
rect -319 238 -307 272
rect -365 232 -307 238
rect -173 272 -115 278
rect -173 238 -161 272
rect -127 238 -115 272
rect -173 232 -115 238
rect 19 272 77 278
rect 19 238 31 272
rect 65 238 77 272
rect 19 232 77 238
rect 211 272 269 278
rect 211 238 223 272
rect 257 238 269 272
rect 211 232 269 238
rect 403 272 461 278
rect 403 238 415 272
rect 449 238 461 272
rect 403 232 461 238
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect -461 -238 -403 -232
rect -461 -272 -449 -238
rect -415 -272 -403 -238
rect -461 -278 -403 -272
rect -269 -238 -211 -232
rect -269 -272 -257 -238
rect -223 -272 -211 -238
rect -269 -278 -211 -272
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -31 -272 -19 -238
rect -77 -278 -19 -272
rect 115 -238 173 -232
rect 115 -272 127 -238
rect 161 -272 173 -238
rect 115 -278 173 -272
rect 307 -238 365 -232
rect 307 -272 319 -238
rect 353 -272 365 -238
rect 307 -278 365 -272
rect -461 -346 -403 -340
rect -461 -380 -449 -346
rect -415 -380 -403 -346
rect -461 -386 -403 -380
rect -269 -346 -211 -340
rect -269 -380 -257 -346
rect -223 -380 -211 -346
rect -269 -386 -211 -380
rect -77 -346 -19 -340
rect -77 -380 -65 -346
rect -31 -380 -19 -346
rect -77 -386 -19 -380
rect 115 -346 173 -340
rect 115 -380 127 -346
rect 161 -380 173 -346
rect 115 -386 173 -380
rect 307 -346 365 -340
rect 307 -380 319 -346
rect 353 -380 365 -346
rect 307 -386 365 -380
rect -503 -430 -457 -418
rect -503 -806 -497 -430
rect -463 -806 -457 -430
rect -503 -818 -457 -806
rect -407 -430 -361 -418
rect -407 -806 -401 -430
rect -367 -806 -361 -430
rect -407 -818 -361 -806
rect -311 -430 -265 -418
rect -311 -806 -305 -430
rect -271 -806 -265 -430
rect -311 -818 -265 -806
rect -215 -430 -169 -418
rect -215 -806 -209 -430
rect -175 -806 -169 -430
rect -215 -818 -169 -806
rect -119 -430 -73 -418
rect -119 -806 -113 -430
rect -79 -806 -73 -430
rect -119 -818 -73 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 73 -430 119 -418
rect 73 -806 79 -430
rect 113 -806 119 -430
rect 73 -818 119 -806
rect 169 -430 215 -418
rect 169 -806 175 -430
rect 209 -806 215 -430
rect 169 -818 215 -806
rect 265 -430 311 -418
rect 265 -806 271 -430
rect 305 -806 311 -430
rect 265 -818 311 -806
rect 361 -430 407 -418
rect 361 -806 367 -430
rect 401 -806 407 -430
rect 361 -818 407 -806
rect 457 -430 503 -418
rect 457 -806 463 -430
rect 497 -806 503 -430
rect 457 -818 503 -806
rect -365 -856 -307 -850
rect -365 -890 -353 -856
rect -319 -890 -307 -856
rect -365 -896 -307 -890
rect -173 -856 -115 -850
rect -173 -890 -161 -856
rect -127 -890 -115 -856
rect -173 -896 -115 -890
rect 19 -856 77 -850
rect 19 -890 31 -856
rect 65 -890 77 -856
rect 19 -896 77 -890
rect 211 -856 269 -850
rect 211 -890 223 -856
rect 257 -890 269 -856
rect 211 -896 269 -890
rect 403 -856 461 -850
rect 403 -890 415 -856
rect 449 -890 461 -856
rect 403 -896 461 -890
rect -365 -964 -307 -958
rect -365 -998 -353 -964
rect -319 -998 -307 -964
rect -365 -1004 -307 -998
rect -173 -964 -115 -958
rect -173 -998 -161 -964
rect -127 -998 -115 -964
rect -173 -1004 -115 -998
rect 19 -964 77 -958
rect 19 -998 31 -964
rect 65 -998 77 -964
rect 19 -1004 77 -998
rect 211 -964 269 -958
rect 211 -998 223 -964
rect 257 -998 269 -964
rect 211 -1004 269 -998
rect 403 -964 461 -958
rect 403 -998 415 -964
rect 449 -998 461 -964
rect 403 -1004 461 -998
rect -503 -1048 -457 -1036
rect -503 -1424 -497 -1048
rect -463 -1424 -457 -1048
rect -503 -1436 -457 -1424
rect -407 -1048 -361 -1036
rect -407 -1424 -401 -1048
rect -367 -1424 -361 -1048
rect -407 -1436 -361 -1424
rect -311 -1048 -265 -1036
rect -311 -1424 -305 -1048
rect -271 -1424 -265 -1048
rect -311 -1436 -265 -1424
rect -215 -1048 -169 -1036
rect -215 -1424 -209 -1048
rect -175 -1424 -169 -1048
rect -215 -1436 -169 -1424
rect -119 -1048 -73 -1036
rect -119 -1424 -113 -1048
rect -79 -1424 -73 -1048
rect -119 -1436 -73 -1424
rect -23 -1048 23 -1036
rect -23 -1424 -17 -1048
rect 17 -1424 23 -1048
rect -23 -1436 23 -1424
rect 73 -1048 119 -1036
rect 73 -1424 79 -1048
rect 113 -1424 119 -1048
rect 73 -1436 119 -1424
rect 169 -1048 215 -1036
rect 169 -1424 175 -1048
rect 209 -1424 215 -1048
rect 169 -1436 215 -1424
rect 265 -1048 311 -1036
rect 265 -1424 271 -1048
rect 305 -1424 311 -1048
rect 265 -1436 311 -1424
rect 361 -1048 407 -1036
rect 361 -1424 367 -1048
rect 401 -1424 407 -1048
rect 361 -1436 407 -1424
rect 457 -1048 503 -1036
rect 457 -1424 463 -1048
rect 497 -1424 503 -1048
rect 457 -1436 503 -1424
rect -461 -1474 -403 -1468
rect -461 -1508 -449 -1474
rect -415 -1508 -403 -1474
rect -461 -1514 -403 -1508
rect -269 -1474 -211 -1468
rect -269 -1508 -257 -1474
rect -223 -1508 -211 -1474
rect -269 -1514 -211 -1508
rect -77 -1474 -19 -1468
rect -77 -1508 -65 -1474
rect -31 -1508 -19 -1474
rect -77 -1514 -19 -1508
rect 115 -1474 173 -1468
rect 115 -1508 127 -1474
rect 161 -1508 173 -1474
rect 115 -1514 173 -1508
rect 307 -1474 365 -1468
rect 307 -1508 319 -1474
rect 353 -1508 365 -1474
rect 307 -1514 365 -1508
<< properties >>
string FIXED_BBOX -594 -1593 594 1593
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 5 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
