* SPICE3 file created from eigth_mirror.ext - technology: sky130A

X0 mirror_p_0/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1 m3_100_0# I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2 m3_100_0# I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3 mirror_p_0/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4 mirror_p_0/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5 mirror_p_0/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6 m3_100_0# I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7 m3_100_0# I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8 m3_100_0# I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9 mirror_p_0/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10 mirror_p_0/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11 m3_100_0# I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12 mirror_p_0/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13 m3_100_0# I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14 mirror_p_0/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15 m3_100_0# I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X16 mirror_p_0/m1_n92_1078# I_In I_In m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X17 I_In I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X18 mirror_p_0/m1_n92_1078# I_In I_In m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X19 I_In I_In mirror_p_0/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X20 mirror_p_1/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X21 m3_100_0# I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X22 m3_100_0# I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X23 mirror_p_1/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X24 mirror_p_1/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X25 mirror_p_1/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X26 m3_100_0# I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X27 m3_100_0# I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X28 m3_100_0# I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X29 mirror_p_1/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X30 mirror_p_1/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X31 m3_100_0# I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X32 mirror_p_1/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X33 m3_100_0# I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X34 mirror_p_1/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X35 m3_100_0# I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X36 mirror_p_1/m1_n92_1078# I_In I_out_0 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X37 I_out_0 I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X38 mirror_p_1/m1_n92_1078# I_In I_out_0 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X39 I_out_0 I_In mirror_p_1/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X40 mirror_p_2/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X41 m3_100_0# I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X42 m3_100_0# I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X43 mirror_p_2/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X44 mirror_p_2/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X45 mirror_p_2/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X46 m3_100_0# I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X47 m3_100_0# I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X48 m3_100_0# I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X49 mirror_p_2/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X50 mirror_p_2/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X51 m3_100_0# I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X52 mirror_p_2/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X53 m3_100_0# I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X54 mirror_p_2/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X55 m3_100_0# I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X56 mirror_p_2/m1_n92_1078# I_In I_out_1 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X57 I_out_1 I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X58 mirror_p_2/m1_n92_1078# I_In I_out_1 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X59 I_out_1 I_In mirror_p_2/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X60 mirror_p_3/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X61 m3_100_0# I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X62 m3_100_0# I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X63 mirror_p_3/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X64 mirror_p_3/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X65 mirror_p_3/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X66 m3_100_0# I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X67 m3_100_0# I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X68 m3_100_0# I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X69 mirror_p_3/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X70 mirror_p_3/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X71 m3_100_0# I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X72 mirror_p_3/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X73 m3_100_0# I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X74 mirror_p_3/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X75 m3_100_0# I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X76 mirror_p_3/m1_n92_1078# I_In I_out_2 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X77 I_out_2 I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X78 mirror_p_3/m1_n92_1078# I_In I_out_2 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X79 I_out_2 I_In mirror_p_3/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X80 mirror_p_4/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X81 m3_100_0# I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X82 m3_100_0# I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X83 mirror_p_4/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X84 mirror_p_4/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X85 mirror_p_4/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X86 m3_100_0# I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X87 m3_100_0# I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X88 m3_100_0# I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X89 mirror_p_4/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X90 mirror_p_4/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X91 m3_100_0# I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X92 mirror_p_4/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X93 m3_100_0# I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X94 mirror_p_4/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X95 m3_100_0# I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X96 mirror_p_4/m1_n92_1078# I_In I_out_3 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X97 I_out_3 I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X98 mirror_p_4/m1_n92_1078# I_In I_out_3 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X99 I_out_3 I_In mirror_p_4/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X100 mirror_p_6/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X101 m3_100_0# I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X102 m3_100_0# I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X103 mirror_p_6/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X104 mirror_p_6/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X105 mirror_p_6/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X106 m3_100_0# I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X107 m3_100_0# I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X108 m3_100_0# I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X109 mirror_p_6/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X110 mirror_p_6/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X111 m3_100_0# I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X112 mirror_p_6/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X113 m3_100_0# I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X114 mirror_p_6/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X115 m3_100_0# I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X116 mirror_p_6/m1_n92_1078# I_In I_out_7 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X117 I_out_7 I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X118 mirror_p_6/m1_n92_1078# I_In I_out_7 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X119 I_out_7 I_In mirror_p_6/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X120 mirror_p_7/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X121 m3_100_0# I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X122 m3_100_0# I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X123 mirror_p_7/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X124 mirror_p_7/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X125 mirror_p_7/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X126 m3_100_0# I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X127 m3_100_0# I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X128 m3_100_0# I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X129 mirror_p_7/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X130 mirror_p_7/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X131 m3_100_0# I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X132 mirror_p_7/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X133 m3_100_0# I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X134 mirror_p_7/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X135 m3_100_0# I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X136 mirror_p_7/m1_n92_1078# I_In I_out_6 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X137 I_out_6 I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X138 mirror_p_7/m1_n92_1078# I_In I_out_6 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X139 I_out_6 I_In mirror_p_7/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X140 mirror_p_8/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X141 m3_100_0# I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X142 m3_100_0# I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X143 mirror_p_8/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X144 mirror_p_8/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X145 mirror_p_8/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X146 m3_100_0# I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X147 m3_100_0# I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X148 m3_100_0# I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X149 mirror_p_8/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X150 mirror_p_8/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X151 m3_100_0# I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X152 mirror_p_8/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X153 m3_100_0# I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X154 mirror_p_8/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X155 m3_100_0# I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X156 mirror_p_8/m1_n92_1078# I_In I_out_5 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X157 I_out_5 I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X158 mirror_p_8/m1_n92_1078# I_In I_out_5 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X159 I_out_5 I_In mirror_p_8/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X160 mirror_p_9/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X161 m3_100_0# I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X162 m3_100_0# I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X163 mirror_p_9/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X164 mirror_p_9/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X165 mirror_p_9/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X166 m3_100_0# I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X167 m3_100_0# I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X168 m3_100_0# I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X169 mirror_p_9/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X170 mirror_p_9/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X171 m3_100_0# I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X172 mirror_p_9/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X173 m3_100_0# I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X174 mirror_p_9/m1_n92_1078# I_In m3_100_0# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X175 m3_100_0# I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X176 mirror_p_9/m1_n92_1078# I_In I_out_4 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X177 I_out_4 I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X178 mirror_p_9/m1_n92_1078# I_In I_out_4 m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
X179 I_out_4 I_In mirror_p_9/m1_n92_1078# m3_100_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=200000u
