magic
tech sky130B
magscale 1 2
timestamp 1654072472
<< error_s >>
rect 117 642 175 648
rect 235 642 293 648
rect 353 642 411 648
rect 471 642 529 648
rect 589 642 647 648
rect 707 642 765 648
rect 825 642 883 648
rect 943 642 1001 648
rect 1061 642 1119 648
rect 1179 642 1237 648
rect 1297 642 1355 648
rect 1415 642 1473 648
rect 117 608 129 642
rect 235 608 247 642
rect 353 608 365 642
rect 471 608 483 642
rect 589 608 601 642
rect 707 608 719 642
rect 825 608 837 642
rect 943 608 955 642
rect 1061 608 1073 642
rect 1179 608 1191 642
rect 1297 608 1309 642
rect 1415 608 1427 642
rect 117 602 175 608
rect 235 602 293 608
rect 353 602 411 608
rect 471 602 529 608
rect 589 602 647 608
rect 707 602 765 608
rect 825 602 883 608
rect 943 602 1001 608
rect 1061 602 1119 608
rect 1179 602 1237 608
rect 1297 602 1355 608
rect 1415 602 1473 608
rect 117 132 175 138
rect 235 132 293 138
rect 353 132 411 138
rect 471 132 529 138
rect 589 132 647 138
rect 707 132 765 138
rect 825 132 883 138
rect 943 132 1001 138
rect 1061 132 1119 138
rect 1179 132 1237 138
rect 1297 132 1355 138
rect 1415 132 1473 138
rect 117 98 129 132
rect 235 98 247 132
rect 353 98 365 132
rect 471 98 483 132
rect 589 98 601 132
rect 707 98 719 132
rect 825 98 837 132
rect 943 98 955 132
rect 1061 98 1073 132
rect 1179 98 1191 132
rect 1297 98 1309 132
rect 1415 98 1427 132
rect 117 92 175 98
rect 235 92 293 98
rect 353 92 411 98
rect 471 92 529 98
rect 589 92 647 98
rect 707 92 765 98
rect 825 92 883 98
rect 943 92 1001 98
rect 1061 92 1119 98
rect 1179 92 1237 98
rect 1297 92 1355 98
rect 1415 92 1473 98
<< metal1 >>
rect 168 410 178 570
rect 232 410 242 570
rect 404 410 414 570
rect 468 410 478 570
rect 640 410 650 570
rect 704 410 714 570
rect 876 410 886 570
rect 940 410 950 570
rect 1112 410 1122 570
rect 1176 410 1186 570
rect 1348 410 1358 570
rect 1412 410 1422 570
rect 50 170 60 330
rect 114 170 124 330
rect 286 170 296 330
rect 350 170 360 330
rect 522 170 532 330
rect 586 170 596 330
rect 758 170 768 330
rect 822 170 832 330
rect 994 170 1004 330
rect 1058 170 1068 330
rect 1230 170 1240 330
rect 1294 170 1304 330
rect 1466 170 1476 330
rect 1530 170 1540 330
<< via1 >>
rect 178 410 232 570
rect 414 410 468 570
rect 650 410 704 570
rect 886 410 940 570
rect 1122 410 1176 570
rect 1358 410 1412 570
rect 60 170 114 330
rect 296 170 350 330
rect 532 170 586 330
rect 768 170 822 330
rect 1004 170 1058 330
rect 1240 170 1294 330
rect 1476 170 1530 330
<< metal2 >>
rect 178 570 232 580
rect 178 400 232 410
rect 414 570 468 580
rect 414 400 468 410
rect 650 570 704 580
rect 650 400 704 410
rect 886 570 940 580
rect 886 400 940 410
rect 1122 570 1176 580
rect 1122 400 1176 410
rect 1358 570 1412 580
rect 1358 400 1412 410
rect 60 330 114 340
rect 60 160 114 170
rect 296 330 350 340
rect 296 160 350 170
rect 532 330 586 340
rect 532 160 586 170
rect 768 330 822 340
rect 768 160 822 170
rect 1004 330 1058 340
rect 1004 160 1058 170
rect 1240 330 1294 340
rect 1240 160 1294 170
rect 1476 330 1530 340
rect 1476 160 1530 170
use sky130_fd_pr__nfet_01v8_lvt_HR8DH9  sky130_fd_pr__nfet_01v8_lvt_HR8DH9_0
timestamp 1654072472
transform 1 0 795 0 1 370
box -875 -410 875 410
<< end >>
