magic
tech sky130A
magscale 1 2
timestamp 1645802395
<< metal3 >>
rect -1350 1272 1349 1300
rect -1350 -1272 1265 1272
rect 1329 -1272 1349 1272
rect -1350 -1300 1349 -1272
<< via3 >>
rect 1265 -1272 1329 1272
<< mimcap >>
rect -1250 1160 1150 1200
rect -1250 -1160 -1210 1160
rect 1110 -1160 1150 1160
rect -1250 -1200 1150 -1160
<< mimcapcontact >>
rect -1210 -1160 1110 1160
<< metal4 >>
rect 1249 1272 1345 1288
rect -1211 1160 1111 1161
rect -1211 -1160 -1210 1160
rect 1110 -1160 1111 1160
rect -1211 -1161 1111 -1160
rect 1249 -1272 1265 1272
rect 1329 -1272 1345 1272
rect 1249 -1288 1345 -1272
<< properties >>
string FIXED_BBOX -1350 -1300 1250 1300
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 12 l 12 val 297.12 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
