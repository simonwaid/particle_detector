magic
tech sky130A
magscale 1 2
timestamp 1647868710
<< locali >>
rect 240 1150 1480 1200
rect 1440 650 1480 1150
rect 1590 750 1600 1200
rect 2190 920 2320 1030
rect 1590 740 2300 750
rect 1440 250 1600 650
rect 1440 160 1630 250
rect 1440 110 1710 160
rect 1440 40 1600 110
<< viali >>
rect 1630 160 1770 250
<< metal1 >>
rect 360 1060 1840 1120
rect 330 800 340 1000
rect 400 800 410 1000
rect 530 800 540 1000
rect 600 800 610 1000
rect 720 800 730 1000
rect 790 800 800 1000
rect 910 800 920 1000
rect 980 800 990 1000
rect 1110 800 1120 1000
rect 1180 800 1190 1000
rect 1310 800 1320 1000
rect 1380 800 1390 1000
rect 1500 860 1580 1060
rect 1660 900 1670 1030
rect 1730 900 1740 1030
rect 1500 800 1800 860
rect 420 230 430 430
rect 490 230 500 430
rect 620 230 630 430
rect 690 230 700 430
rect 820 230 830 430
rect 890 230 900 430
rect 1010 230 1020 430
rect 1080 230 1090 430
rect 1210 230 1220 430
rect 1280 230 1290 430
rect 1500 160 1580 800
rect 1740 530 1750 600
rect 1900 530 1910 600
rect 1630 350 1640 480
rect 1700 350 1710 480
rect 1770 320 1830 530
rect 360 100 1580 160
rect 1618 250 1782 256
rect 1618 160 1630 250
rect 1770 160 1782 250
rect 1618 154 1782 160
<< via1 >>
rect 340 800 400 1000
rect 540 800 600 1000
rect 730 800 790 1000
rect 920 800 980 1000
rect 1120 800 1180 1000
rect 1320 800 1380 1000
rect 1670 900 1730 1030
rect 430 230 490 430
rect 630 230 690 430
rect 830 230 890 430
rect 1020 230 1080 430
rect 1220 230 1280 430
rect 1750 530 1900 600
rect 1640 350 1700 480
rect 1630 160 1770 250
<< metal2 >>
rect 1670 1030 1730 1040
rect 340 1000 400 1010
rect 540 1000 600 1010
rect 730 1000 790 1010
rect 920 1000 980 1010
rect 1120 1000 1180 1010
rect 1320 1000 1380 1010
rect 1520 1000 1670 1030
rect 400 800 540 1000
rect 600 800 730 1000
rect 790 800 920 1000
rect 980 800 1120 1000
rect 1180 800 1320 1000
rect 1380 920 1670 1000
rect 1380 800 1630 920
rect 1730 920 1750 1030
rect 1670 890 1730 900
rect 340 790 400 800
rect 540 790 600 800
rect 730 790 790 800
rect 920 790 980 800
rect 1120 790 1180 800
rect 1320 790 1380 800
rect 1520 610 1630 800
rect 1520 600 1900 610
rect 1520 530 1750 600
rect 1750 520 1900 530
rect 1640 480 1700 490
rect 430 430 490 440
rect 630 430 690 440
rect 830 430 890 440
rect 1020 430 1080 440
rect 1220 430 1280 440
rect 350 230 430 430
rect 490 230 630 430
rect 690 230 830 430
rect 890 230 1020 430
rect 1080 230 1220 430
rect 1280 350 1640 430
rect 1700 350 1710 430
rect 1280 260 1710 350
rect 1280 250 1770 260
rect 1280 230 1630 250
rect 430 220 490 230
rect 630 220 690 230
rect 830 220 890 230
rect 1020 220 1080 230
rect 1220 220 1280 230
rect 1630 150 1770 160
use sky130_fd_pr__nfet_01v8_U3V43Z  sky130_fd_pr__nfet_01v8_U3V43Z_0
timestamp 1647868710
transform 1 0 1936 0 1 440
box -396 -260 396 260
use sky130_fd_pr__nfet_01v8_lvt_E9U3PA  sky130_fd_pr__nfet_01v8_lvt_E9U3PA_0
timestamp 1647868710
transform 1 0 857 0 1 610
box -657 -610 657 610
use sky130_fd_pr__pfet_01v8_QDYTZD  sky130_fd_pr__pfet_01v8_QDYTZD_1
timestamp 1647868710
transform 1 0 1956 0 1 969
box -396 -269 396 269
<< end >>
