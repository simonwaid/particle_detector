magic
tech sky130B
magscale 1 2
timestamp 1654683408
<< nwell >>
rect 230 1916 3080 1982
rect 248 1902 278 1916
rect 440 1902 470 1916
rect 632 1902 662 1916
rect 824 1902 854 1916
rect 1016 1902 1046 1916
rect 1208 1902 1238 1916
rect 1400 1902 1430 1916
rect 1592 1910 1622 1916
rect 1784 1910 1814 1916
rect 1976 1910 2006 1916
rect 2168 1910 2198 1916
rect 2360 1910 2390 1916
rect 2552 1910 2582 1916
rect 2744 1910 2774 1916
rect 2936 1910 2966 1916
rect 344 1454 374 1466
rect 536 1454 566 1466
rect 728 1454 758 1466
rect 920 1454 950 1464
rect 1112 1454 1142 1466
rect 1304 1454 1334 1464
rect 1496 1454 1526 1464
rect 1688 1454 1718 1466
rect 1880 1454 1910 1466
rect 2072 1454 2102 1468
rect 2264 1454 2294 1468
rect 2456 1454 2486 1466
rect 2648 1454 2678 1466
rect 2840 1454 2870 1464
rect 3032 1454 3062 1466
rect 230 1388 3080 1454
rect 230 1280 3080 1346
rect 344 1268 374 1280
rect 536 1268 566 1280
rect 728 1268 758 1280
rect 920 1270 950 1280
rect 1112 1268 1142 1280
rect 1304 1270 1334 1280
rect 1496 1270 1526 1280
rect 1688 1268 1718 1280
rect 1880 1268 1910 1280
rect 2072 1266 2102 1280
rect 2264 1266 2294 1280
rect 2456 1268 2486 1280
rect 2648 1268 2678 1280
rect 2840 1270 2870 1280
rect 3032 1268 3062 1280
rect 248 818 278 832
rect 440 818 470 832
rect 632 818 662 832
rect 824 818 854 832
rect 1016 818 1046 832
rect 1208 818 1238 832
rect 1400 818 1430 832
rect 1592 818 1622 824
rect 1784 818 1814 824
rect 1976 818 2006 824
rect 2168 818 2198 824
rect 2360 818 2390 824
rect 2552 818 2582 824
rect 2744 818 2774 824
rect 2936 818 2966 824
rect 230 752 3080 818
rect 230 644 3080 710
rect 248 630 278 644
rect 440 630 470 644
rect 632 630 662 644
rect 824 630 854 644
rect 1016 630 1046 644
rect 1208 630 1238 644
rect 1400 630 1430 644
rect 1592 638 1622 644
rect 1784 638 1814 644
rect 1976 638 2006 644
rect 2168 638 2198 644
rect 2360 638 2390 644
rect 2552 638 2582 644
rect 2744 638 2774 644
rect 2936 638 2966 644
rect 344 182 374 194
rect 536 182 566 194
rect 728 182 758 194
rect 920 182 950 192
rect 1112 182 1142 194
rect 1304 182 1334 192
rect 1496 182 1526 192
rect 1688 182 1718 194
rect 1880 182 1910 194
rect 2072 182 2102 196
rect 2264 182 2294 196
rect 2456 182 2486 194
rect 2648 182 2678 194
rect 2840 182 2870 192
rect 3032 182 3062 194
rect 230 116 3080 182
<< poly >>
rect 230 1966 3080 1982
rect 230 1932 246 1966
rect 280 1932 438 1966
rect 472 1932 630 1966
rect 664 1932 822 1966
rect 856 1932 1014 1966
rect 1048 1932 1206 1966
rect 1240 1932 1398 1966
rect 1432 1932 1590 1966
rect 1624 1932 1782 1966
rect 1816 1932 1974 1966
rect 2008 1932 2166 1966
rect 2200 1932 2358 1966
rect 2392 1932 2550 1966
rect 2584 1932 2742 1966
rect 2776 1932 2934 1966
rect 2968 1932 3080 1966
rect 230 1916 3080 1932
rect 248 1902 278 1916
rect 440 1902 470 1916
rect 632 1902 662 1916
rect 824 1902 854 1916
rect 1016 1902 1046 1916
rect 1208 1902 1238 1916
rect 1400 1902 1430 1916
rect 1592 1910 1622 1916
rect 1784 1910 1814 1916
rect 1976 1910 2006 1916
rect 2168 1910 2198 1916
rect 2360 1910 2390 1916
rect 2552 1910 2582 1916
rect 2744 1910 2774 1916
rect 2936 1910 2966 1916
rect 344 1454 374 1466
rect 536 1454 566 1466
rect 728 1454 758 1466
rect 920 1454 950 1464
rect 1112 1454 1142 1466
rect 1304 1454 1334 1464
rect 1496 1454 1526 1464
rect 1688 1454 1718 1466
rect 1880 1454 1910 1466
rect 2072 1454 2102 1468
rect 2264 1454 2294 1468
rect 2456 1454 2486 1466
rect 2648 1454 2678 1466
rect 2840 1454 2870 1464
rect 3032 1454 3062 1466
rect 230 1438 3080 1454
rect 230 1404 342 1438
rect 376 1404 534 1438
rect 568 1404 726 1438
rect 760 1404 918 1438
rect 952 1404 1110 1438
rect 1144 1404 1302 1438
rect 1336 1404 1494 1438
rect 1528 1404 1686 1438
rect 1720 1404 1878 1438
rect 1912 1404 2070 1438
rect 2104 1404 2262 1438
rect 2296 1404 2454 1438
rect 2488 1404 2646 1438
rect 2680 1404 2838 1438
rect 2872 1404 3030 1438
rect 3064 1404 3080 1438
rect 230 1388 3080 1404
rect 230 1330 3080 1346
rect 230 1296 342 1330
rect 376 1296 534 1330
rect 568 1296 726 1330
rect 760 1296 918 1330
rect 952 1296 1110 1330
rect 1144 1296 1302 1330
rect 1336 1296 1494 1330
rect 1528 1296 1686 1330
rect 1720 1296 1878 1330
rect 1912 1296 2070 1330
rect 2104 1296 2262 1330
rect 2296 1296 2454 1330
rect 2488 1296 2646 1330
rect 2680 1296 2838 1330
rect 2872 1296 3030 1330
rect 3064 1296 3080 1330
rect 230 1280 3080 1296
rect 344 1268 374 1280
rect 536 1268 566 1280
rect 728 1268 758 1280
rect 920 1270 950 1280
rect 1112 1268 1142 1280
rect 1304 1270 1334 1280
rect 1496 1270 1526 1280
rect 1688 1268 1718 1280
rect 1880 1268 1910 1280
rect 2072 1266 2102 1280
rect 2264 1266 2294 1280
rect 2456 1268 2486 1280
rect 2648 1268 2678 1280
rect 2840 1270 2870 1280
rect 3032 1268 3062 1280
rect 248 818 278 832
rect 440 818 470 832
rect 632 818 662 832
rect 824 818 854 832
rect 1016 818 1046 832
rect 1208 818 1238 832
rect 1400 818 1430 832
rect 1592 818 1622 824
rect 1784 818 1814 824
rect 1976 818 2006 824
rect 2168 818 2198 824
rect 2360 818 2390 824
rect 2552 818 2582 824
rect 2744 818 2774 824
rect 2936 818 2966 824
rect 230 802 3080 818
rect 230 768 246 802
rect 280 768 438 802
rect 472 768 630 802
rect 664 768 822 802
rect 856 768 1014 802
rect 1048 768 1206 802
rect 1240 768 1398 802
rect 1432 768 1590 802
rect 1624 768 1782 802
rect 1816 768 1974 802
rect 2008 768 2166 802
rect 2200 768 2358 802
rect 2392 768 2550 802
rect 2584 768 2742 802
rect 2776 768 2934 802
rect 2968 768 3080 802
rect 230 752 3080 768
rect 230 694 3080 710
rect 230 660 246 694
rect 280 660 438 694
rect 472 660 630 694
rect 664 660 822 694
rect 856 660 1014 694
rect 1048 660 1206 694
rect 1240 660 1398 694
rect 1432 660 1590 694
rect 1624 660 1782 694
rect 1816 660 1974 694
rect 2008 660 2166 694
rect 2200 660 2358 694
rect 2392 660 2550 694
rect 2584 660 2742 694
rect 2776 660 2934 694
rect 2968 660 3080 694
rect 230 644 3080 660
rect 248 630 278 644
rect 440 630 470 644
rect 632 630 662 644
rect 824 630 854 644
rect 1016 630 1046 644
rect 1208 630 1238 644
rect 1400 630 1430 644
rect 1592 638 1622 644
rect 1784 638 1814 644
rect 1976 638 2006 644
rect 2168 638 2198 644
rect 2360 638 2390 644
rect 2552 638 2582 644
rect 2744 638 2774 644
rect 2936 638 2966 644
rect 344 182 374 194
rect 536 182 566 194
rect 728 182 758 194
rect 920 182 950 192
rect 1112 182 1142 194
rect 1304 182 1334 192
rect 1496 182 1526 192
rect 1688 182 1718 194
rect 1880 182 1910 194
rect 2072 182 2102 196
rect 2264 182 2294 196
rect 2456 182 2486 194
rect 2648 182 2678 194
rect 2840 182 2870 192
rect 3032 182 3062 194
rect 230 166 3080 182
rect 230 132 342 166
rect 376 132 534 166
rect 568 132 726 166
rect 760 132 918 166
rect 952 132 1110 166
rect 1144 132 1302 166
rect 1336 132 1494 166
rect 1528 132 1686 166
rect 1720 132 1878 166
rect 1912 132 2070 166
rect 2104 132 2262 166
rect 2296 132 2454 166
rect 2488 132 2646 166
rect 2680 132 2838 166
rect 2872 132 3030 166
rect 3064 132 3080 166
rect 230 116 3080 132
<< polycont >>
rect 246 1932 280 1966
rect 438 1932 472 1966
rect 630 1932 664 1966
rect 822 1932 856 1966
rect 1014 1932 1048 1966
rect 1206 1932 1240 1966
rect 1398 1932 1432 1966
rect 1590 1932 1624 1966
rect 1782 1932 1816 1966
rect 1974 1932 2008 1966
rect 2166 1932 2200 1966
rect 2358 1932 2392 1966
rect 2550 1932 2584 1966
rect 2742 1932 2776 1966
rect 2934 1932 2968 1966
rect 342 1404 376 1438
rect 534 1404 568 1438
rect 726 1404 760 1438
rect 918 1404 952 1438
rect 1110 1404 1144 1438
rect 1302 1404 1336 1438
rect 1494 1404 1528 1438
rect 1686 1404 1720 1438
rect 1878 1404 1912 1438
rect 2070 1404 2104 1438
rect 2262 1404 2296 1438
rect 2454 1404 2488 1438
rect 2646 1404 2680 1438
rect 2838 1404 2872 1438
rect 3030 1404 3064 1438
rect 342 1296 376 1330
rect 534 1296 568 1330
rect 726 1296 760 1330
rect 918 1296 952 1330
rect 1110 1296 1144 1330
rect 1302 1296 1336 1330
rect 1494 1296 1528 1330
rect 1686 1296 1720 1330
rect 1878 1296 1912 1330
rect 2070 1296 2104 1330
rect 2262 1296 2296 1330
rect 2454 1296 2488 1330
rect 2646 1296 2680 1330
rect 2838 1296 2872 1330
rect 3030 1296 3064 1330
rect 246 768 280 802
rect 438 768 472 802
rect 630 768 664 802
rect 822 768 856 802
rect 1014 768 1048 802
rect 1206 768 1240 802
rect 1398 768 1432 802
rect 1590 768 1624 802
rect 1782 768 1816 802
rect 1974 768 2008 802
rect 2166 768 2200 802
rect 2358 768 2392 802
rect 2550 768 2584 802
rect 2742 768 2776 802
rect 2934 768 2968 802
rect 246 660 280 694
rect 438 660 472 694
rect 630 660 664 694
rect 822 660 856 694
rect 1014 660 1048 694
rect 1206 660 1240 694
rect 1398 660 1432 694
rect 1590 660 1624 694
rect 1782 660 1816 694
rect 1974 660 2008 694
rect 2166 660 2200 694
rect 2358 660 2392 694
rect 2550 660 2584 694
rect 2742 660 2776 694
rect 2934 660 2968 694
rect 342 132 376 166
rect 534 132 568 166
rect 726 132 760 166
rect 918 132 952 166
rect 1110 132 1144 166
rect 1302 132 1336 166
rect 1494 132 1528 166
rect 1686 132 1720 166
rect 1878 132 1912 166
rect 2070 132 2104 166
rect 2262 132 2296 166
rect 2454 132 2488 166
rect 2646 132 2680 166
rect 2838 132 2872 166
rect 3030 132 3064 166
<< locali >>
rect 230 1932 246 1966
rect 280 1932 438 1966
rect 472 1932 630 1966
rect 664 1932 822 1966
rect 856 1932 1014 1966
rect 1048 1932 1206 1966
rect 1240 1932 1398 1966
rect 1432 1932 1590 1966
rect 1624 1932 1782 1966
rect 1816 1932 1974 1966
rect 2008 1932 2166 1966
rect 2200 1932 2358 1966
rect 2392 1932 2550 1966
rect 2584 1932 2742 1966
rect 2776 1932 2934 1966
rect 2968 1932 3080 1966
rect 230 1404 342 1438
rect 376 1404 534 1438
rect 568 1404 726 1438
rect 760 1404 918 1438
rect 952 1404 1110 1438
rect 1144 1404 1302 1438
rect 1336 1404 1494 1438
rect 1528 1404 1686 1438
rect 1720 1404 1878 1438
rect 1912 1404 2070 1438
rect 2104 1404 2262 1438
rect 2296 1404 2454 1438
rect 2488 1404 2646 1438
rect 2680 1404 2838 1438
rect 2872 1404 3030 1438
rect 3064 1404 3080 1438
rect 230 1296 342 1330
rect 376 1296 534 1330
rect 568 1296 726 1330
rect 760 1296 918 1330
rect 952 1296 1110 1330
rect 1144 1296 1302 1330
rect 1336 1296 1494 1330
rect 1528 1296 1686 1330
rect 1720 1296 1878 1330
rect 1912 1296 2070 1330
rect 2104 1296 2262 1330
rect 2296 1296 2454 1330
rect 2488 1296 2646 1330
rect 2680 1296 2838 1330
rect 2872 1296 3030 1330
rect 3064 1296 3080 1330
rect 230 768 246 802
rect 280 768 438 802
rect 472 768 630 802
rect 664 768 822 802
rect 856 768 1014 802
rect 1048 768 1206 802
rect 1240 768 1398 802
rect 1432 768 1590 802
rect 1624 768 1782 802
rect 1816 768 1974 802
rect 2008 768 2166 802
rect 2200 768 2358 802
rect 2392 768 2550 802
rect 2584 768 2742 802
rect 2776 768 2934 802
rect 2968 768 3080 802
rect 230 660 246 694
rect 280 660 438 694
rect 472 660 630 694
rect 664 660 822 694
rect 856 660 1014 694
rect 1048 660 1206 694
rect 1240 660 1398 694
rect 1432 660 1590 694
rect 1624 660 1782 694
rect 1816 660 1974 694
rect 2008 660 2166 694
rect 2200 660 2358 694
rect 2392 660 2550 694
rect 2584 660 2742 694
rect 2776 660 2934 694
rect 2968 660 3080 694
rect 230 132 342 166
rect 376 132 534 166
rect 568 132 726 166
rect 760 132 918 166
rect 952 132 1110 166
rect 1144 132 1302 166
rect 1336 132 1494 166
rect 1528 132 1686 166
rect 1720 132 1878 166
rect 1912 132 2070 166
rect 2104 132 2262 166
rect 2296 132 2454 166
rect 2488 132 2646 166
rect 2680 132 2838 166
rect 2872 132 3030 166
rect 3064 132 3080 166
<< viali >>
rect 246 1932 280 1966
rect 438 1932 472 1966
rect 630 1932 664 1966
rect 822 1932 856 1966
rect 1014 1932 1048 1966
rect 1206 1932 1240 1966
rect 1398 1932 1432 1966
rect 1590 1932 1624 1966
rect 1782 1932 1816 1966
rect 1974 1932 2008 1966
rect 2166 1932 2200 1966
rect 2358 1932 2392 1966
rect 2550 1932 2584 1966
rect 2742 1932 2776 1966
rect 2934 1932 2968 1966
rect 342 1404 376 1438
rect 534 1404 568 1438
rect 726 1404 760 1438
rect 918 1404 952 1438
rect 1110 1404 1144 1438
rect 1302 1404 1336 1438
rect 1494 1404 1528 1438
rect 1686 1404 1720 1438
rect 1878 1404 1912 1438
rect 2070 1404 2104 1438
rect 2262 1404 2296 1438
rect 2454 1404 2488 1438
rect 2646 1404 2680 1438
rect 2838 1404 2872 1438
rect 3030 1404 3064 1438
rect 342 1296 376 1330
rect 534 1296 568 1330
rect 726 1296 760 1330
rect 918 1296 952 1330
rect 1110 1296 1144 1330
rect 1302 1296 1336 1330
rect 1494 1296 1528 1330
rect 1686 1296 1720 1330
rect 1878 1296 1912 1330
rect 2070 1296 2104 1330
rect 2262 1296 2296 1330
rect 2454 1296 2488 1330
rect 2646 1296 2680 1330
rect 2838 1296 2872 1330
rect 3030 1296 3064 1330
rect 246 768 280 802
rect 438 768 472 802
rect 630 768 664 802
rect 822 768 856 802
rect 1014 768 1048 802
rect 1206 768 1240 802
rect 1398 768 1432 802
rect 1590 768 1624 802
rect 1782 768 1816 802
rect 1974 768 2008 802
rect 2166 768 2200 802
rect 2358 768 2392 802
rect 2550 768 2584 802
rect 2742 768 2776 802
rect 2934 768 2968 802
rect 246 660 280 694
rect 438 660 472 694
rect 630 660 664 694
rect 822 660 856 694
rect 1014 660 1048 694
rect 1206 660 1240 694
rect 1398 660 1432 694
rect 1590 660 1624 694
rect 1782 660 1816 694
rect 1974 660 2008 694
rect 2166 660 2200 694
rect 2358 660 2392 694
rect 2550 660 2584 694
rect 2742 660 2776 694
rect 2934 660 2968 694
rect 342 132 376 166
rect 534 132 568 166
rect 726 132 760 166
rect 918 132 952 166
rect 1110 132 1144 166
rect 1302 132 1336 166
rect 1494 132 1528 166
rect 1686 132 1720 166
rect 1878 132 1912 166
rect 2070 132 2104 166
rect 2262 132 2296 166
rect 2454 132 2488 166
rect 2646 132 2680 166
rect 2838 132 2872 166
rect 3030 132 3064 166
<< metal1 >>
rect 110 1966 3200 2020
rect 110 1932 246 1966
rect 280 1932 438 1966
rect 472 1932 630 1966
rect 664 1932 822 1966
rect 856 1932 1014 1966
rect 1048 1932 1206 1966
rect 1240 1932 1398 1966
rect 1432 1932 1590 1966
rect 1624 1932 1782 1966
rect 1816 1932 1974 1966
rect 2008 1932 2166 1966
rect 2200 1932 2358 1966
rect 2392 1932 2550 1966
rect 2584 1932 2742 1966
rect 2776 1932 2934 1966
rect 2968 1932 3200 1966
rect 110 1920 3200 1932
rect 274 1710 284 1886
rect 338 1710 348 1886
rect 466 1710 476 1886
rect 530 1710 540 1886
rect 658 1710 668 1886
rect 722 1710 732 1886
rect 850 1710 860 1886
rect 914 1710 924 1886
rect 1042 1710 1052 1886
rect 1106 1710 1116 1886
rect 1234 1710 1244 1886
rect 1298 1710 1308 1886
rect 1426 1710 1436 1886
rect 1490 1710 1500 1886
rect 1618 1710 1628 1886
rect 1682 1710 1692 1886
rect 1810 1710 1820 1886
rect 1874 1710 1884 1886
rect 2002 1710 2012 1886
rect 2066 1710 2076 1886
rect 2194 1710 2204 1886
rect 2258 1710 2268 1886
rect 2386 1710 2396 1886
rect 2450 1710 2460 1886
rect 2578 1710 2588 1886
rect 2642 1710 2652 1886
rect 2770 1710 2780 1886
rect 2834 1710 2844 1886
rect 2962 1710 2972 1886
rect 3026 1710 3036 1886
rect 178 1484 188 1660
rect 242 1484 252 1660
rect 370 1484 380 1660
rect 434 1484 444 1660
rect 562 1484 572 1660
rect 626 1484 636 1660
rect 754 1484 764 1660
rect 818 1484 828 1660
rect 946 1484 956 1660
rect 1010 1484 1020 1660
rect 1138 1484 1148 1660
rect 1202 1484 1212 1660
rect 1330 1484 1340 1660
rect 1394 1484 1404 1660
rect 1522 1484 1532 1660
rect 1586 1484 1596 1660
rect 1714 1484 1724 1660
rect 1778 1484 1788 1660
rect 1906 1484 1916 1660
rect 1970 1484 1980 1660
rect 2098 1484 2108 1660
rect 2162 1484 2172 1660
rect 2290 1484 2300 1660
rect 2354 1484 2364 1660
rect 2482 1484 2492 1660
rect 2546 1484 2556 1660
rect 2674 1484 2684 1660
rect 2738 1484 2748 1660
rect 2866 1484 2876 1660
rect 2930 1484 2940 1660
rect 3058 1484 3068 1660
rect 3122 1484 3132 1660
rect 110 1438 3200 1450
rect 110 1404 342 1438
rect 376 1404 534 1438
rect 568 1404 726 1438
rect 760 1404 918 1438
rect 952 1404 1110 1438
rect 1144 1404 1302 1438
rect 1336 1404 1494 1438
rect 1528 1404 1686 1438
rect 1720 1404 1878 1438
rect 1912 1404 2070 1438
rect 2104 1404 2262 1438
rect 2296 1404 2454 1438
rect 2488 1404 2646 1438
rect 2680 1404 2838 1438
rect 2872 1404 3030 1438
rect 3064 1404 3200 1438
rect 110 1330 3200 1404
rect 110 1296 342 1330
rect 376 1296 534 1330
rect 568 1296 726 1330
rect 760 1296 918 1330
rect 952 1296 1110 1330
rect 1144 1296 1302 1330
rect 1336 1296 1494 1330
rect 1528 1296 1686 1330
rect 1720 1296 1878 1330
rect 1912 1296 2070 1330
rect 2104 1296 2262 1330
rect 2296 1296 2454 1330
rect 2488 1296 2646 1330
rect 2680 1296 2838 1330
rect 2872 1296 3030 1330
rect 3064 1296 3200 1330
rect 110 1290 3200 1296
rect 178 1074 188 1250
rect 242 1074 252 1250
rect 370 1074 380 1250
rect 434 1074 444 1250
rect 562 1074 572 1250
rect 626 1074 636 1250
rect 754 1074 764 1250
rect 818 1074 828 1250
rect 946 1074 956 1250
rect 1010 1074 1020 1250
rect 1138 1074 1148 1250
rect 1202 1074 1212 1250
rect 1330 1074 1340 1250
rect 1394 1074 1404 1250
rect 1522 1074 1532 1250
rect 1586 1074 1596 1250
rect 1714 1074 1724 1250
rect 1778 1074 1788 1250
rect 1906 1074 1916 1250
rect 1970 1074 1980 1250
rect 2098 1074 2108 1250
rect 2162 1074 2172 1250
rect 2290 1074 2300 1250
rect 2354 1074 2364 1250
rect 2482 1074 2492 1250
rect 2546 1074 2556 1250
rect 2674 1074 2684 1250
rect 2738 1074 2748 1250
rect 2866 1074 2876 1250
rect 2930 1074 2940 1250
rect 3058 1074 3068 1250
rect 3122 1074 3132 1250
rect 274 848 284 1024
rect 338 848 348 1024
rect 466 848 476 1024
rect 530 848 540 1024
rect 658 848 668 1024
rect 722 848 732 1024
rect 850 848 860 1024
rect 914 848 924 1024
rect 1042 848 1052 1024
rect 1106 848 1116 1024
rect 1234 848 1244 1024
rect 1298 848 1308 1024
rect 1426 848 1436 1024
rect 1490 848 1500 1024
rect 1618 848 1628 1024
rect 1682 848 1692 1024
rect 1810 848 1820 1024
rect 1874 848 1884 1024
rect 2002 848 2012 1024
rect 2066 848 2076 1024
rect 2194 848 2204 1024
rect 2258 848 2268 1024
rect 2386 848 2396 1024
rect 2450 848 2460 1024
rect 2578 848 2588 1024
rect 2642 848 2652 1024
rect 2770 848 2780 1024
rect 2834 848 2844 1024
rect 2962 848 2972 1024
rect 3026 848 3036 1024
rect 110 802 3200 810
rect 110 768 246 802
rect 280 768 438 802
rect 472 768 630 802
rect 664 768 822 802
rect 856 768 1014 802
rect 1048 768 1206 802
rect 1240 768 1398 802
rect 1432 768 1590 802
rect 1624 768 1782 802
rect 1816 768 1974 802
rect 2008 768 2166 802
rect 2200 768 2358 802
rect 2392 768 2550 802
rect 2584 768 2742 802
rect 2776 768 2934 802
rect 2968 768 3200 802
rect 110 694 3200 768
rect 110 660 246 694
rect 280 660 438 694
rect 472 660 630 694
rect 664 660 822 694
rect 856 660 1014 694
rect 1048 660 1206 694
rect 1240 660 1398 694
rect 1432 660 1590 694
rect 1624 660 1782 694
rect 1816 660 1974 694
rect 2008 660 2166 694
rect 2200 660 2358 694
rect 2392 660 2550 694
rect 2584 660 2742 694
rect 2776 660 2934 694
rect 2968 660 3200 694
rect 110 650 3200 660
rect 274 438 284 614
rect 338 438 348 614
rect 466 438 476 614
rect 530 438 540 614
rect 658 438 668 614
rect 722 438 732 614
rect 850 438 860 614
rect 914 438 924 614
rect 1042 438 1052 614
rect 1106 438 1116 614
rect 1234 438 1244 614
rect 1298 438 1308 614
rect 1426 438 1436 614
rect 1490 438 1500 614
rect 1618 438 1628 614
rect 1682 438 1692 614
rect 1810 438 1820 614
rect 1874 438 1884 614
rect 2002 438 2012 614
rect 2066 438 2076 614
rect 2194 438 2204 614
rect 2258 438 2268 614
rect 2386 438 2396 614
rect 2450 438 2460 614
rect 2578 438 2588 614
rect 2642 438 2652 614
rect 2770 438 2780 614
rect 2834 438 2844 614
rect 2962 438 2972 614
rect 3026 438 3036 614
rect 178 212 188 388
rect 242 212 252 388
rect 370 212 380 388
rect 434 212 444 388
rect 562 212 572 388
rect 626 212 636 388
rect 754 212 764 388
rect 818 212 828 388
rect 946 212 956 388
rect 1010 212 1020 388
rect 1138 212 1148 388
rect 1202 212 1212 388
rect 1330 212 1340 388
rect 1394 212 1404 388
rect 1522 212 1532 388
rect 1586 212 1596 388
rect 1714 212 1724 388
rect 1778 212 1788 388
rect 1906 212 1916 388
rect 1970 212 1980 388
rect 2098 212 2108 388
rect 2162 212 2172 388
rect 2290 212 2300 388
rect 2354 212 2364 388
rect 2482 212 2492 388
rect 2546 212 2556 388
rect 2674 212 2684 388
rect 2738 212 2748 388
rect 2866 212 2876 388
rect 2930 212 2940 388
rect 3058 212 3068 388
rect 3122 212 3132 388
rect 110 166 3200 180
rect 110 132 342 166
rect 376 132 534 166
rect 568 132 726 166
rect 760 132 918 166
rect 952 132 1110 166
rect 1144 132 1302 166
rect 1336 132 1494 166
rect 1528 132 1686 166
rect 1720 132 1878 166
rect 1912 132 2070 166
rect 2104 132 2262 166
rect 2296 132 2454 166
rect 2488 132 2646 166
rect 2680 132 2838 166
rect 2872 132 3030 166
rect 3064 132 3200 166
rect 110 80 3200 132
<< via1 >>
rect 284 1710 338 1886
rect 476 1710 530 1886
rect 668 1710 722 1886
rect 860 1710 914 1886
rect 1052 1710 1106 1886
rect 1244 1710 1298 1886
rect 1436 1710 1490 1886
rect 1628 1710 1682 1886
rect 1820 1710 1874 1886
rect 2012 1710 2066 1886
rect 2204 1710 2258 1886
rect 2396 1710 2450 1886
rect 2588 1710 2642 1886
rect 2780 1710 2834 1886
rect 2972 1710 3026 1886
rect 188 1484 242 1660
rect 380 1484 434 1660
rect 572 1484 626 1660
rect 764 1484 818 1660
rect 956 1484 1010 1660
rect 1148 1484 1202 1660
rect 1340 1484 1394 1660
rect 1532 1484 1586 1660
rect 1724 1484 1778 1660
rect 1916 1484 1970 1660
rect 2108 1484 2162 1660
rect 2300 1484 2354 1660
rect 2492 1484 2546 1660
rect 2684 1484 2738 1660
rect 2876 1484 2930 1660
rect 3068 1484 3122 1660
rect 188 1074 242 1250
rect 380 1074 434 1250
rect 572 1074 626 1250
rect 764 1074 818 1250
rect 956 1074 1010 1250
rect 1148 1074 1202 1250
rect 1340 1074 1394 1250
rect 1532 1074 1586 1250
rect 1724 1074 1778 1250
rect 1916 1074 1970 1250
rect 2108 1074 2162 1250
rect 2300 1074 2354 1250
rect 2492 1074 2546 1250
rect 2684 1074 2738 1250
rect 2876 1074 2930 1250
rect 3068 1074 3122 1250
rect 284 848 338 1024
rect 476 848 530 1024
rect 668 848 722 1024
rect 860 848 914 1024
rect 1052 848 1106 1024
rect 1244 848 1298 1024
rect 1436 848 1490 1024
rect 1628 848 1682 1024
rect 1820 848 1874 1024
rect 2012 848 2066 1024
rect 2204 848 2258 1024
rect 2396 848 2450 1024
rect 2588 848 2642 1024
rect 2780 848 2834 1024
rect 2972 848 3026 1024
rect 284 438 338 614
rect 476 438 530 614
rect 668 438 722 614
rect 860 438 914 614
rect 1052 438 1106 614
rect 1244 438 1298 614
rect 1436 438 1490 614
rect 1628 438 1682 614
rect 1820 438 1874 614
rect 2012 438 2066 614
rect 2204 438 2258 614
rect 2396 438 2450 614
rect 2588 438 2642 614
rect 2780 438 2834 614
rect 2972 438 3026 614
rect 188 212 242 388
rect 380 212 434 388
rect 572 212 626 388
rect 764 212 818 388
rect 956 212 1010 388
rect 1148 212 1202 388
rect 1340 212 1394 388
rect 1532 212 1586 388
rect 1724 212 1778 388
rect 1916 212 1970 388
rect 2108 212 2162 388
rect 2300 212 2354 388
rect 2492 212 2546 388
rect 2684 212 2738 388
rect 2876 212 2930 388
rect 3068 212 3122 388
<< metal2 >>
rect 284 1886 3026 1896
rect 338 1736 476 1886
rect 284 1700 338 1710
rect 530 1736 668 1886
rect 476 1700 530 1710
rect 722 1736 860 1886
rect 668 1700 722 1710
rect 914 1736 1052 1886
rect 860 1700 914 1710
rect 1106 1736 1244 1886
rect 1052 1700 1106 1710
rect 1298 1736 1436 1886
rect 1244 1700 1298 1710
rect 1490 1736 1628 1886
rect 1436 1700 1490 1710
rect 1682 1736 1820 1886
rect 1628 1700 1682 1710
rect 1874 1736 2012 1886
rect 1820 1700 1874 1710
rect 2066 1736 2204 1886
rect 2012 1700 2066 1710
rect 2258 1736 2396 1886
rect 2204 1700 2258 1710
rect 2450 1736 2588 1886
rect 2396 1700 2450 1710
rect 2642 1736 2780 1886
rect 2588 1700 2642 1710
rect 2834 1736 2972 1886
rect 2780 1700 2834 1710
rect 2972 1700 3026 1710
rect 188 1660 242 1670
rect 380 1660 434 1670
rect 242 1484 380 1634
rect 572 1660 626 1670
rect 434 1484 572 1634
rect 764 1660 818 1670
rect 626 1484 764 1634
rect 956 1660 1010 1670
rect 818 1484 956 1634
rect 1148 1660 1202 1670
rect 1010 1484 1148 1634
rect 1340 1660 1394 1670
rect 1202 1484 1340 1634
rect 1532 1660 1586 1670
rect 1394 1484 1532 1634
rect 1724 1660 1778 1670
rect 1586 1484 1724 1634
rect 1916 1660 1970 1670
rect 1778 1484 1916 1634
rect 2108 1660 2162 1670
rect 1970 1484 2108 1634
rect 2300 1660 2354 1670
rect 2162 1484 2300 1634
rect 2492 1660 2546 1670
rect 2354 1484 2492 1634
rect 2684 1660 2738 1670
rect 2546 1484 2684 1634
rect 2876 1660 2930 1670
rect 2738 1484 2876 1634
rect 3068 1660 3122 1670
rect 2930 1484 3068 1634
rect 188 1474 3122 1484
rect 188 1250 3122 1260
rect 242 1100 380 1250
rect 188 1064 242 1074
rect 434 1100 572 1250
rect 380 1064 434 1074
rect 626 1100 764 1250
rect 572 1064 626 1074
rect 818 1100 956 1250
rect 764 1064 818 1074
rect 1010 1100 1148 1250
rect 956 1064 1010 1074
rect 1202 1100 1340 1250
rect 1148 1064 1202 1074
rect 1394 1100 1532 1250
rect 1340 1064 1394 1074
rect 1586 1100 1724 1250
rect 1532 1064 1586 1074
rect 1778 1100 1916 1250
rect 1724 1064 1778 1074
rect 1970 1100 2108 1250
rect 1916 1064 1970 1074
rect 2162 1100 2300 1250
rect 2108 1064 2162 1074
rect 2354 1100 2492 1250
rect 2300 1064 2354 1074
rect 2546 1100 2684 1250
rect 2492 1064 2546 1074
rect 2738 1100 2876 1250
rect 2684 1064 2738 1074
rect 2930 1100 3068 1250
rect 2876 1064 2930 1074
rect 3068 1064 3122 1074
rect 284 1024 338 1034
rect 476 1024 530 1034
rect 338 848 476 998
rect 668 1024 722 1034
rect 530 848 668 998
rect 860 1024 914 1034
rect 722 848 860 998
rect 1052 1024 1106 1034
rect 914 848 1052 998
rect 1244 1024 1298 1034
rect 1106 848 1244 998
rect 1436 1024 1490 1034
rect 1298 848 1436 998
rect 1628 1024 1682 1034
rect 1490 848 1628 998
rect 1820 1024 1874 1034
rect 1682 848 1820 998
rect 2012 1024 2066 1034
rect 1874 848 2012 998
rect 2204 1024 2258 1034
rect 2066 848 2204 998
rect 2396 1024 2450 1034
rect 2258 848 2396 998
rect 2588 1024 2642 1034
rect 2450 848 2588 998
rect 2780 1024 2834 1034
rect 2642 848 2780 998
rect 2972 1024 3026 1034
rect 2834 848 2972 998
rect 284 838 3026 848
rect 284 614 3026 624
rect 338 464 476 614
rect 284 428 338 438
rect 530 464 668 614
rect 476 428 530 438
rect 722 464 860 614
rect 668 428 722 438
rect 914 464 1052 614
rect 860 428 914 438
rect 1106 464 1244 614
rect 1052 428 1106 438
rect 1298 464 1436 614
rect 1244 428 1298 438
rect 1490 464 1628 614
rect 1436 428 1490 438
rect 1682 464 1820 614
rect 1628 428 1682 438
rect 1874 464 2012 614
rect 1820 428 1874 438
rect 2066 464 2204 614
rect 2012 428 2066 438
rect 2258 464 2396 614
rect 2204 428 2258 438
rect 2450 464 2588 614
rect 2396 428 2450 438
rect 2642 464 2780 614
rect 2588 428 2642 438
rect 2834 464 2972 614
rect 2780 428 2834 438
rect 2972 428 3026 438
rect 188 388 242 398
rect 380 388 434 398
rect 242 212 380 362
rect 572 388 626 398
rect 434 212 572 362
rect 764 388 818 398
rect 626 212 764 362
rect 956 388 1010 398
rect 818 212 956 362
rect 1148 388 1202 398
rect 1010 212 1148 362
rect 1340 388 1394 398
rect 1202 212 1340 362
rect 1532 388 1586 398
rect 1394 212 1532 362
rect 1724 388 1778 398
rect 1586 212 1724 362
rect 1916 388 1970 398
rect 1778 212 1916 362
rect 2108 388 2162 398
rect 1970 212 2108 362
rect 2300 388 2354 398
rect 2162 212 2300 362
rect 2492 388 2546 398
rect 2354 212 2492 362
rect 2684 388 2738 398
rect 2546 212 2684 362
rect 2876 388 2930 398
rect 2738 212 2876 362
rect 3068 388 3122 398
rect 2930 212 3068 362
rect 188 202 3122 212
use sky130_fd_pr__pfet_01v8_VCB4SW  sky130_fd_pr__pfet_01v8_VCB4SW_0
timestamp 1654683408
transform 1 0 1655 0 1 1049
box -1607 -1055 1607 1055
<< end >>
