magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< error_p >>
rect -1181 1199 -1123 1205
rect -989 1199 -931 1205
rect -797 1199 -739 1205
rect -605 1199 -547 1205
rect -413 1199 -355 1205
rect -221 1199 -163 1205
rect -29 1199 29 1205
rect 163 1199 221 1205
rect 355 1199 413 1205
rect 547 1199 605 1205
rect 739 1199 797 1205
rect 931 1199 989 1205
rect 1123 1199 1181 1205
rect -1181 1165 -1169 1199
rect -989 1165 -977 1199
rect -797 1165 -785 1199
rect -605 1165 -593 1199
rect -413 1165 -401 1199
rect -221 1165 -209 1199
rect -29 1165 -17 1199
rect 163 1165 175 1199
rect 355 1165 367 1199
rect 547 1165 559 1199
rect 739 1165 751 1199
rect 931 1165 943 1199
rect 1123 1165 1135 1199
rect -1181 1159 -1123 1165
rect -989 1159 -931 1165
rect -797 1159 -739 1165
rect -605 1159 -547 1165
rect -413 1159 -355 1165
rect -221 1159 -163 1165
rect -29 1159 29 1165
rect 163 1159 221 1165
rect 355 1159 413 1165
rect 547 1159 605 1165
rect 739 1159 797 1165
rect 931 1159 989 1165
rect 1123 1159 1181 1165
rect -1085 689 -1027 695
rect -893 689 -835 695
rect -701 689 -643 695
rect -509 689 -451 695
rect -317 689 -259 695
rect -125 689 -67 695
rect 67 689 125 695
rect 259 689 317 695
rect 451 689 509 695
rect 643 689 701 695
rect 835 689 893 695
rect 1027 689 1085 695
rect -1085 655 -1073 689
rect -893 655 -881 689
rect -701 655 -689 689
rect -509 655 -497 689
rect -317 655 -305 689
rect -125 655 -113 689
rect 67 655 79 689
rect 259 655 271 689
rect 451 655 463 689
rect 643 655 655 689
rect 835 655 847 689
rect 1027 655 1039 689
rect -1085 649 -1027 655
rect -893 649 -835 655
rect -701 649 -643 655
rect -509 649 -451 655
rect -317 649 -259 655
rect -125 649 -67 655
rect 67 649 125 655
rect 259 649 317 655
rect 451 649 509 655
rect 643 649 701 655
rect 835 649 893 655
rect 1027 649 1085 655
rect -1085 581 -1027 587
rect -893 581 -835 587
rect -701 581 -643 587
rect -509 581 -451 587
rect -317 581 -259 587
rect -125 581 -67 587
rect 67 581 125 587
rect 259 581 317 587
rect 451 581 509 587
rect 643 581 701 587
rect 835 581 893 587
rect 1027 581 1085 587
rect -1085 547 -1073 581
rect -893 547 -881 581
rect -701 547 -689 581
rect -509 547 -497 581
rect -317 547 -305 581
rect -125 547 -113 581
rect 67 547 79 581
rect 259 547 271 581
rect 451 547 463 581
rect 643 547 655 581
rect 835 547 847 581
rect 1027 547 1039 581
rect -1085 541 -1027 547
rect -893 541 -835 547
rect -701 541 -643 547
rect -509 541 -451 547
rect -317 541 -259 547
rect -125 541 -67 547
rect 67 541 125 547
rect 259 541 317 547
rect 451 541 509 547
rect 643 541 701 547
rect 835 541 893 547
rect 1027 541 1085 547
rect -1181 71 -1123 77
rect -989 71 -931 77
rect -797 71 -739 77
rect -605 71 -547 77
rect -413 71 -355 77
rect -221 71 -163 77
rect -29 71 29 77
rect 163 71 221 77
rect 355 71 413 77
rect 547 71 605 77
rect 739 71 797 77
rect 931 71 989 77
rect 1123 71 1181 77
rect -1181 37 -1169 71
rect -989 37 -977 71
rect -797 37 -785 71
rect -605 37 -593 71
rect -413 37 -401 71
rect -221 37 -209 71
rect -29 37 -17 71
rect 163 37 175 71
rect 355 37 367 71
rect 547 37 559 71
rect 739 37 751 71
rect 931 37 943 71
rect 1123 37 1135 71
rect -1181 31 -1123 37
rect -989 31 -931 37
rect -797 31 -739 37
rect -605 31 -547 37
rect -413 31 -355 37
rect -221 31 -163 37
rect -29 31 29 37
rect 163 31 221 37
rect 355 31 413 37
rect 547 31 605 37
rect 739 31 797 37
rect 931 31 989 37
rect 1123 31 1181 37
rect -1181 -37 -1123 -31
rect -989 -37 -931 -31
rect -797 -37 -739 -31
rect -605 -37 -547 -31
rect -413 -37 -355 -31
rect -221 -37 -163 -31
rect -29 -37 29 -31
rect 163 -37 221 -31
rect 355 -37 413 -31
rect 547 -37 605 -31
rect 739 -37 797 -31
rect 931 -37 989 -31
rect 1123 -37 1181 -31
rect -1181 -71 -1169 -37
rect -989 -71 -977 -37
rect -797 -71 -785 -37
rect -605 -71 -593 -37
rect -413 -71 -401 -37
rect -221 -71 -209 -37
rect -29 -71 -17 -37
rect 163 -71 175 -37
rect 355 -71 367 -37
rect 547 -71 559 -37
rect 739 -71 751 -37
rect 931 -71 943 -37
rect 1123 -71 1135 -37
rect -1181 -77 -1123 -71
rect -989 -77 -931 -71
rect -797 -77 -739 -71
rect -605 -77 -547 -71
rect -413 -77 -355 -71
rect -221 -77 -163 -71
rect -29 -77 29 -71
rect 163 -77 221 -71
rect 355 -77 413 -71
rect 547 -77 605 -71
rect 739 -77 797 -71
rect 931 -77 989 -71
rect 1123 -77 1181 -71
rect -1085 -547 -1027 -541
rect -893 -547 -835 -541
rect -701 -547 -643 -541
rect -509 -547 -451 -541
rect -317 -547 -259 -541
rect -125 -547 -67 -541
rect 67 -547 125 -541
rect 259 -547 317 -541
rect 451 -547 509 -541
rect 643 -547 701 -541
rect 835 -547 893 -541
rect 1027 -547 1085 -541
rect -1085 -581 -1073 -547
rect -893 -581 -881 -547
rect -701 -581 -689 -547
rect -509 -581 -497 -547
rect -317 -581 -305 -547
rect -125 -581 -113 -547
rect 67 -581 79 -547
rect 259 -581 271 -547
rect 451 -581 463 -547
rect 643 -581 655 -547
rect 835 -581 847 -547
rect 1027 -581 1039 -547
rect -1085 -587 -1027 -581
rect -893 -587 -835 -581
rect -701 -587 -643 -581
rect -509 -587 -451 -581
rect -317 -587 -259 -581
rect -125 -587 -67 -581
rect 67 -587 125 -581
rect 259 -587 317 -581
rect 451 -587 509 -581
rect 643 -587 701 -581
rect 835 -587 893 -581
rect 1027 -587 1085 -581
rect -1085 -655 -1027 -649
rect -893 -655 -835 -649
rect -701 -655 -643 -649
rect -509 -655 -451 -649
rect -317 -655 -259 -649
rect -125 -655 -67 -649
rect 67 -655 125 -649
rect 259 -655 317 -649
rect 451 -655 509 -649
rect 643 -655 701 -649
rect 835 -655 893 -649
rect 1027 -655 1085 -649
rect -1085 -689 -1073 -655
rect -893 -689 -881 -655
rect -701 -689 -689 -655
rect -509 -689 -497 -655
rect -317 -689 -305 -655
rect -125 -689 -113 -655
rect 67 -689 79 -655
rect 259 -689 271 -655
rect 451 -689 463 -655
rect 643 -689 655 -655
rect 835 -689 847 -655
rect 1027 -689 1039 -655
rect -1085 -695 -1027 -689
rect -893 -695 -835 -689
rect -701 -695 -643 -689
rect -509 -695 -451 -689
rect -317 -695 -259 -689
rect -125 -695 -67 -689
rect 67 -695 125 -689
rect 259 -695 317 -689
rect 451 -695 509 -689
rect 643 -695 701 -689
rect 835 -695 893 -689
rect 1027 -695 1085 -689
rect -1181 -1165 -1123 -1159
rect -989 -1165 -931 -1159
rect -797 -1165 -739 -1159
rect -605 -1165 -547 -1159
rect -413 -1165 -355 -1159
rect -221 -1165 -163 -1159
rect -29 -1165 29 -1159
rect 163 -1165 221 -1159
rect 355 -1165 413 -1159
rect 547 -1165 605 -1159
rect 739 -1165 797 -1159
rect 931 -1165 989 -1159
rect 1123 -1165 1181 -1159
rect -1181 -1199 -1169 -1165
rect -989 -1199 -977 -1165
rect -797 -1199 -785 -1165
rect -605 -1199 -593 -1165
rect -413 -1199 -401 -1165
rect -221 -1199 -209 -1165
rect -29 -1199 -17 -1165
rect 163 -1199 175 -1165
rect 355 -1199 367 -1165
rect 547 -1199 559 -1165
rect 739 -1199 751 -1165
rect 931 -1199 943 -1165
rect 1123 -1199 1135 -1165
rect -1181 -1205 -1123 -1199
rect -989 -1205 -931 -1199
rect -797 -1205 -739 -1199
rect -605 -1205 -547 -1199
rect -413 -1205 -355 -1199
rect -221 -1205 -163 -1199
rect -29 -1205 29 -1199
rect 163 -1205 221 -1199
rect 355 -1205 413 -1199
rect 547 -1205 605 -1199
rect 739 -1205 797 -1199
rect 931 -1205 989 -1199
rect 1123 -1205 1181 -1199
<< nmos >>
rect -1167 727 -1137 1127
rect -1071 727 -1041 1127
rect -975 727 -945 1127
rect -879 727 -849 1127
rect -783 727 -753 1127
rect -687 727 -657 1127
rect -591 727 -561 1127
rect -495 727 -465 1127
rect -399 727 -369 1127
rect -303 727 -273 1127
rect -207 727 -177 1127
rect -111 727 -81 1127
rect -15 727 15 1127
rect 81 727 111 1127
rect 177 727 207 1127
rect 273 727 303 1127
rect 369 727 399 1127
rect 465 727 495 1127
rect 561 727 591 1127
rect 657 727 687 1127
rect 753 727 783 1127
rect 849 727 879 1127
rect 945 727 975 1127
rect 1041 727 1071 1127
rect 1137 727 1167 1127
rect -1167 109 -1137 509
rect -1071 109 -1041 509
rect -975 109 -945 509
rect -879 109 -849 509
rect -783 109 -753 509
rect -687 109 -657 509
rect -591 109 -561 509
rect -495 109 -465 509
rect -399 109 -369 509
rect -303 109 -273 509
rect -207 109 -177 509
rect -111 109 -81 509
rect -15 109 15 509
rect 81 109 111 509
rect 177 109 207 509
rect 273 109 303 509
rect 369 109 399 509
rect 465 109 495 509
rect 561 109 591 509
rect 657 109 687 509
rect 753 109 783 509
rect 849 109 879 509
rect 945 109 975 509
rect 1041 109 1071 509
rect 1137 109 1167 509
rect -1167 -509 -1137 -109
rect -1071 -509 -1041 -109
rect -975 -509 -945 -109
rect -879 -509 -849 -109
rect -783 -509 -753 -109
rect -687 -509 -657 -109
rect -591 -509 -561 -109
rect -495 -509 -465 -109
rect -399 -509 -369 -109
rect -303 -509 -273 -109
rect -207 -509 -177 -109
rect -111 -509 -81 -109
rect -15 -509 15 -109
rect 81 -509 111 -109
rect 177 -509 207 -109
rect 273 -509 303 -109
rect 369 -509 399 -109
rect 465 -509 495 -109
rect 561 -509 591 -109
rect 657 -509 687 -109
rect 753 -509 783 -109
rect 849 -509 879 -109
rect 945 -509 975 -109
rect 1041 -509 1071 -109
rect 1137 -509 1167 -109
rect -1167 -1127 -1137 -727
rect -1071 -1127 -1041 -727
rect -975 -1127 -945 -727
rect -879 -1127 -849 -727
rect -783 -1127 -753 -727
rect -687 -1127 -657 -727
rect -591 -1127 -561 -727
rect -495 -1127 -465 -727
rect -399 -1127 -369 -727
rect -303 -1127 -273 -727
rect -207 -1127 -177 -727
rect -111 -1127 -81 -727
rect -15 -1127 15 -727
rect 81 -1127 111 -727
rect 177 -1127 207 -727
rect 273 -1127 303 -727
rect 369 -1127 399 -727
rect 465 -1127 495 -727
rect 561 -1127 591 -727
rect 657 -1127 687 -727
rect 753 -1127 783 -727
rect 849 -1127 879 -727
rect 945 -1127 975 -727
rect 1041 -1127 1071 -727
rect 1137 -1127 1167 -727
<< ndiff >>
rect -1229 1115 -1167 1127
rect -1229 739 -1217 1115
rect -1183 739 -1167 1115
rect -1229 727 -1167 739
rect -1137 1115 -1071 1127
rect -1137 739 -1121 1115
rect -1087 739 -1071 1115
rect -1137 727 -1071 739
rect -1041 1115 -975 1127
rect -1041 739 -1025 1115
rect -991 739 -975 1115
rect -1041 727 -975 739
rect -945 1115 -879 1127
rect -945 739 -929 1115
rect -895 739 -879 1115
rect -945 727 -879 739
rect -849 1115 -783 1127
rect -849 739 -833 1115
rect -799 739 -783 1115
rect -849 727 -783 739
rect -753 1115 -687 1127
rect -753 739 -737 1115
rect -703 739 -687 1115
rect -753 727 -687 739
rect -657 1115 -591 1127
rect -657 739 -641 1115
rect -607 739 -591 1115
rect -657 727 -591 739
rect -561 1115 -495 1127
rect -561 739 -545 1115
rect -511 739 -495 1115
rect -561 727 -495 739
rect -465 1115 -399 1127
rect -465 739 -449 1115
rect -415 739 -399 1115
rect -465 727 -399 739
rect -369 1115 -303 1127
rect -369 739 -353 1115
rect -319 739 -303 1115
rect -369 727 -303 739
rect -273 1115 -207 1127
rect -273 739 -257 1115
rect -223 739 -207 1115
rect -273 727 -207 739
rect -177 1115 -111 1127
rect -177 739 -161 1115
rect -127 739 -111 1115
rect -177 727 -111 739
rect -81 1115 -15 1127
rect -81 739 -65 1115
rect -31 739 -15 1115
rect -81 727 -15 739
rect 15 1115 81 1127
rect 15 739 31 1115
rect 65 739 81 1115
rect 15 727 81 739
rect 111 1115 177 1127
rect 111 739 127 1115
rect 161 739 177 1115
rect 111 727 177 739
rect 207 1115 273 1127
rect 207 739 223 1115
rect 257 739 273 1115
rect 207 727 273 739
rect 303 1115 369 1127
rect 303 739 319 1115
rect 353 739 369 1115
rect 303 727 369 739
rect 399 1115 465 1127
rect 399 739 415 1115
rect 449 739 465 1115
rect 399 727 465 739
rect 495 1115 561 1127
rect 495 739 511 1115
rect 545 739 561 1115
rect 495 727 561 739
rect 591 1115 657 1127
rect 591 739 607 1115
rect 641 739 657 1115
rect 591 727 657 739
rect 687 1115 753 1127
rect 687 739 703 1115
rect 737 739 753 1115
rect 687 727 753 739
rect 783 1115 849 1127
rect 783 739 799 1115
rect 833 739 849 1115
rect 783 727 849 739
rect 879 1115 945 1127
rect 879 739 895 1115
rect 929 739 945 1115
rect 879 727 945 739
rect 975 1115 1041 1127
rect 975 739 991 1115
rect 1025 739 1041 1115
rect 975 727 1041 739
rect 1071 1115 1137 1127
rect 1071 739 1087 1115
rect 1121 739 1137 1115
rect 1071 727 1137 739
rect 1167 1115 1229 1127
rect 1167 739 1183 1115
rect 1217 739 1229 1115
rect 1167 727 1229 739
rect -1229 497 -1167 509
rect -1229 121 -1217 497
rect -1183 121 -1167 497
rect -1229 109 -1167 121
rect -1137 497 -1071 509
rect -1137 121 -1121 497
rect -1087 121 -1071 497
rect -1137 109 -1071 121
rect -1041 497 -975 509
rect -1041 121 -1025 497
rect -991 121 -975 497
rect -1041 109 -975 121
rect -945 497 -879 509
rect -945 121 -929 497
rect -895 121 -879 497
rect -945 109 -879 121
rect -849 497 -783 509
rect -849 121 -833 497
rect -799 121 -783 497
rect -849 109 -783 121
rect -753 497 -687 509
rect -753 121 -737 497
rect -703 121 -687 497
rect -753 109 -687 121
rect -657 497 -591 509
rect -657 121 -641 497
rect -607 121 -591 497
rect -657 109 -591 121
rect -561 497 -495 509
rect -561 121 -545 497
rect -511 121 -495 497
rect -561 109 -495 121
rect -465 497 -399 509
rect -465 121 -449 497
rect -415 121 -399 497
rect -465 109 -399 121
rect -369 497 -303 509
rect -369 121 -353 497
rect -319 121 -303 497
rect -369 109 -303 121
rect -273 497 -207 509
rect -273 121 -257 497
rect -223 121 -207 497
rect -273 109 -207 121
rect -177 497 -111 509
rect -177 121 -161 497
rect -127 121 -111 497
rect -177 109 -111 121
rect -81 497 -15 509
rect -81 121 -65 497
rect -31 121 -15 497
rect -81 109 -15 121
rect 15 497 81 509
rect 15 121 31 497
rect 65 121 81 497
rect 15 109 81 121
rect 111 497 177 509
rect 111 121 127 497
rect 161 121 177 497
rect 111 109 177 121
rect 207 497 273 509
rect 207 121 223 497
rect 257 121 273 497
rect 207 109 273 121
rect 303 497 369 509
rect 303 121 319 497
rect 353 121 369 497
rect 303 109 369 121
rect 399 497 465 509
rect 399 121 415 497
rect 449 121 465 497
rect 399 109 465 121
rect 495 497 561 509
rect 495 121 511 497
rect 545 121 561 497
rect 495 109 561 121
rect 591 497 657 509
rect 591 121 607 497
rect 641 121 657 497
rect 591 109 657 121
rect 687 497 753 509
rect 687 121 703 497
rect 737 121 753 497
rect 687 109 753 121
rect 783 497 849 509
rect 783 121 799 497
rect 833 121 849 497
rect 783 109 849 121
rect 879 497 945 509
rect 879 121 895 497
rect 929 121 945 497
rect 879 109 945 121
rect 975 497 1041 509
rect 975 121 991 497
rect 1025 121 1041 497
rect 975 109 1041 121
rect 1071 497 1137 509
rect 1071 121 1087 497
rect 1121 121 1137 497
rect 1071 109 1137 121
rect 1167 497 1229 509
rect 1167 121 1183 497
rect 1217 121 1229 497
rect 1167 109 1229 121
rect -1229 -121 -1167 -109
rect -1229 -497 -1217 -121
rect -1183 -497 -1167 -121
rect -1229 -509 -1167 -497
rect -1137 -121 -1071 -109
rect -1137 -497 -1121 -121
rect -1087 -497 -1071 -121
rect -1137 -509 -1071 -497
rect -1041 -121 -975 -109
rect -1041 -497 -1025 -121
rect -991 -497 -975 -121
rect -1041 -509 -975 -497
rect -945 -121 -879 -109
rect -945 -497 -929 -121
rect -895 -497 -879 -121
rect -945 -509 -879 -497
rect -849 -121 -783 -109
rect -849 -497 -833 -121
rect -799 -497 -783 -121
rect -849 -509 -783 -497
rect -753 -121 -687 -109
rect -753 -497 -737 -121
rect -703 -497 -687 -121
rect -753 -509 -687 -497
rect -657 -121 -591 -109
rect -657 -497 -641 -121
rect -607 -497 -591 -121
rect -657 -509 -591 -497
rect -561 -121 -495 -109
rect -561 -497 -545 -121
rect -511 -497 -495 -121
rect -561 -509 -495 -497
rect -465 -121 -399 -109
rect -465 -497 -449 -121
rect -415 -497 -399 -121
rect -465 -509 -399 -497
rect -369 -121 -303 -109
rect -369 -497 -353 -121
rect -319 -497 -303 -121
rect -369 -509 -303 -497
rect -273 -121 -207 -109
rect -273 -497 -257 -121
rect -223 -497 -207 -121
rect -273 -509 -207 -497
rect -177 -121 -111 -109
rect -177 -497 -161 -121
rect -127 -497 -111 -121
rect -177 -509 -111 -497
rect -81 -121 -15 -109
rect -81 -497 -65 -121
rect -31 -497 -15 -121
rect -81 -509 -15 -497
rect 15 -121 81 -109
rect 15 -497 31 -121
rect 65 -497 81 -121
rect 15 -509 81 -497
rect 111 -121 177 -109
rect 111 -497 127 -121
rect 161 -497 177 -121
rect 111 -509 177 -497
rect 207 -121 273 -109
rect 207 -497 223 -121
rect 257 -497 273 -121
rect 207 -509 273 -497
rect 303 -121 369 -109
rect 303 -497 319 -121
rect 353 -497 369 -121
rect 303 -509 369 -497
rect 399 -121 465 -109
rect 399 -497 415 -121
rect 449 -497 465 -121
rect 399 -509 465 -497
rect 495 -121 561 -109
rect 495 -497 511 -121
rect 545 -497 561 -121
rect 495 -509 561 -497
rect 591 -121 657 -109
rect 591 -497 607 -121
rect 641 -497 657 -121
rect 591 -509 657 -497
rect 687 -121 753 -109
rect 687 -497 703 -121
rect 737 -497 753 -121
rect 687 -509 753 -497
rect 783 -121 849 -109
rect 783 -497 799 -121
rect 833 -497 849 -121
rect 783 -509 849 -497
rect 879 -121 945 -109
rect 879 -497 895 -121
rect 929 -497 945 -121
rect 879 -509 945 -497
rect 975 -121 1041 -109
rect 975 -497 991 -121
rect 1025 -497 1041 -121
rect 975 -509 1041 -497
rect 1071 -121 1137 -109
rect 1071 -497 1087 -121
rect 1121 -497 1137 -121
rect 1071 -509 1137 -497
rect 1167 -121 1229 -109
rect 1167 -497 1183 -121
rect 1217 -497 1229 -121
rect 1167 -509 1229 -497
rect -1229 -739 -1167 -727
rect -1229 -1115 -1217 -739
rect -1183 -1115 -1167 -739
rect -1229 -1127 -1167 -1115
rect -1137 -739 -1071 -727
rect -1137 -1115 -1121 -739
rect -1087 -1115 -1071 -739
rect -1137 -1127 -1071 -1115
rect -1041 -739 -975 -727
rect -1041 -1115 -1025 -739
rect -991 -1115 -975 -739
rect -1041 -1127 -975 -1115
rect -945 -739 -879 -727
rect -945 -1115 -929 -739
rect -895 -1115 -879 -739
rect -945 -1127 -879 -1115
rect -849 -739 -783 -727
rect -849 -1115 -833 -739
rect -799 -1115 -783 -739
rect -849 -1127 -783 -1115
rect -753 -739 -687 -727
rect -753 -1115 -737 -739
rect -703 -1115 -687 -739
rect -753 -1127 -687 -1115
rect -657 -739 -591 -727
rect -657 -1115 -641 -739
rect -607 -1115 -591 -739
rect -657 -1127 -591 -1115
rect -561 -739 -495 -727
rect -561 -1115 -545 -739
rect -511 -1115 -495 -739
rect -561 -1127 -495 -1115
rect -465 -739 -399 -727
rect -465 -1115 -449 -739
rect -415 -1115 -399 -739
rect -465 -1127 -399 -1115
rect -369 -739 -303 -727
rect -369 -1115 -353 -739
rect -319 -1115 -303 -739
rect -369 -1127 -303 -1115
rect -273 -739 -207 -727
rect -273 -1115 -257 -739
rect -223 -1115 -207 -739
rect -273 -1127 -207 -1115
rect -177 -739 -111 -727
rect -177 -1115 -161 -739
rect -127 -1115 -111 -739
rect -177 -1127 -111 -1115
rect -81 -739 -15 -727
rect -81 -1115 -65 -739
rect -31 -1115 -15 -739
rect -81 -1127 -15 -1115
rect 15 -739 81 -727
rect 15 -1115 31 -739
rect 65 -1115 81 -739
rect 15 -1127 81 -1115
rect 111 -739 177 -727
rect 111 -1115 127 -739
rect 161 -1115 177 -739
rect 111 -1127 177 -1115
rect 207 -739 273 -727
rect 207 -1115 223 -739
rect 257 -1115 273 -739
rect 207 -1127 273 -1115
rect 303 -739 369 -727
rect 303 -1115 319 -739
rect 353 -1115 369 -739
rect 303 -1127 369 -1115
rect 399 -739 465 -727
rect 399 -1115 415 -739
rect 449 -1115 465 -739
rect 399 -1127 465 -1115
rect 495 -739 561 -727
rect 495 -1115 511 -739
rect 545 -1115 561 -739
rect 495 -1127 561 -1115
rect 591 -739 657 -727
rect 591 -1115 607 -739
rect 641 -1115 657 -739
rect 591 -1127 657 -1115
rect 687 -739 753 -727
rect 687 -1115 703 -739
rect 737 -1115 753 -739
rect 687 -1127 753 -1115
rect 783 -739 849 -727
rect 783 -1115 799 -739
rect 833 -1115 849 -739
rect 783 -1127 849 -1115
rect 879 -739 945 -727
rect 879 -1115 895 -739
rect 929 -1115 945 -739
rect 879 -1127 945 -1115
rect 975 -739 1041 -727
rect 975 -1115 991 -739
rect 1025 -1115 1041 -739
rect 975 -1127 1041 -1115
rect 1071 -739 1137 -727
rect 1071 -1115 1087 -739
rect 1121 -1115 1137 -739
rect 1071 -1127 1137 -1115
rect 1167 -739 1229 -727
rect 1167 -1115 1183 -739
rect 1217 -1115 1229 -739
rect 1167 -1127 1229 -1115
<< ndiffc >>
rect -1217 739 -1183 1115
rect -1121 739 -1087 1115
rect -1025 739 -991 1115
rect -929 739 -895 1115
rect -833 739 -799 1115
rect -737 739 -703 1115
rect -641 739 -607 1115
rect -545 739 -511 1115
rect -449 739 -415 1115
rect -353 739 -319 1115
rect -257 739 -223 1115
rect -161 739 -127 1115
rect -65 739 -31 1115
rect 31 739 65 1115
rect 127 739 161 1115
rect 223 739 257 1115
rect 319 739 353 1115
rect 415 739 449 1115
rect 511 739 545 1115
rect 607 739 641 1115
rect 703 739 737 1115
rect 799 739 833 1115
rect 895 739 929 1115
rect 991 739 1025 1115
rect 1087 739 1121 1115
rect 1183 739 1217 1115
rect -1217 121 -1183 497
rect -1121 121 -1087 497
rect -1025 121 -991 497
rect -929 121 -895 497
rect -833 121 -799 497
rect -737 121 -703 497
rect -641 121 -607 497
rect -545 121 -511 497
rect -449 121 -415 497
rect -353 121 -319 497
rect -257 121 -223 497
rect -161 121 -127 497
rect -65 121 -31 497
rect 31 121 65 497
rect 127 121 161 497
rect 223 121 257 497
rect 319 121 353 497
rect 415 121 449 497
rect 511 121 545 497
rect 607 121 641 497
rect 703 121 737 497
rect 799 121 833 497
rect 895 121 929 497
rect 991 121 1025 497
rect 1087 121 1121 497
rect 1183 121 1217 497
rect -1217 -497 -1183 -121
rect -1121 -497 -1087 -121
rect -1025 -497 -991 -121
rect -929 -497 -895 -121
rect -833 -497 -799 -121
rect -737 -497 -703 -121
rect -641 -497 -607 -121
rect -545 -497 -511 -121
rect -449 -497 -415 -121
rect -353 -497 -319 -121
rect -257 -497 -223 -121
rect -161 -497 -127 -121
rect -65 -497 -31 -121
rect 31 -497 65 -121
rect 127 -497 161 -121
rect 223 -497 257 -121
rect 319 -497 353 -121
rect 415 -497 449 -121
rect 511 -497 545 -121
rect 607 -497 641 -121
rect 703 -497 737 -121
rect 799 -497 833 -121
rect 895 -497 929 -121
rect 991 -497 1025 -121
rect 1087 -497 1121 -121
rect 1183 -497 1217 -121
rect -1217 -1115 -1183 -739
rect -1121 -1115 -1087 -739
rect -1025 -1115 -991 -739
rect -929 -1115 -895 -739
rect -833 -1115 -799 -739
rect -737 -1115 -703 -739
rect -641 -1115 -607 -739
rect -545 -1115 -511 -739
rect -449 -1115 -415 -739
rect -353 -1115 -319 -739
rect -257 -1115 -223 -739
rect -161 -1115 -127 -739
rect -65 -1115 -31 -739
rect 31 -1115 65 -739
rect 127 -1115 161 -739
rect 223 -1115 257 -739
rect 319 -1115 353 -739
rect 415 -1115 449 -739
rect 511 -1115 545 -739
rect 607 -1115 641 -739
rect 703 -1115 737 -739
rect 799 -1115 833 -739
rect 895 -1115 929 -739
rect 991 -1115 1025 -739
rect 1087 -1115 1121 -739
rect 1183 -1115 1217 -739
<< psubdiff >>
rect -1331 1267 -1235 1301
rect 1235 1267 1331 1301
rect -1331 1205 -1297 1267
rect 1297 1205 1331 1267
rect -1331 -1267 -1297 -1205
rect 1297 -1267 1331 -1205
rect -1331 -1301 -1235 -1267
rect 1235 -1301 1331 -1267
<< psubdiffcont >>
rect -1235 1267 1235 1301
rect -1331 -1205 -1297 1205
rect 1297 -1205 1331 1205
rect -1235 -1301 1235 -1267
<< poly >>
rect -1185 1199 -1119 1215
rect -1185 1165 -1169 1199
rect -1135 1165 -1119 1199
rect -1185 1149 -1119 1165
rect -993 1199 -927 1215
rect -993 1165 -977 1199
rect -943 1165 -927 1199
rect -1167 1127 -1137 1149
rect -1071 1127 -1041 1153
rect -993 1149 -927 1165
rect -801 1199 -735 1215
rect -801 1165 -785 1199
rect -751 1165 -735 1199
rect -975 1127 -945 1149
rect -879 1127 -849 1153
rect -801 1149 -735 1165
rect -609 1199 -543 1215
rect -609 1165 -593 1199
rect -559 1165 -543 1199
rect -783 1127 -753 1149
rect -687 1127 -657 1153
rect -609 1149 -543 1165
rect -417 1199 -351 1215
rect -417 1165 -401 1199
rect -367 1165 -351 1199
rect -591 1127 -561 1149
rect -495 1127 -465 1153
rect -417 1149 -351 1165
rect -225 1199 -159 1215
rect -225 1165 -209 1199
rect -175 1165 -159 1199
rect -399 1127 -369 1149
rect -303 1127 -273 1153
rect -225 1149 -159 1165
rect -33 1199 33 1215
rect -33 1165 -17 1199
rect 17 1165 33 1199
rect -207 1127 -177 1149
rect -111 1127 -81 1153
rect -33 1149 33 1165
rect 159 1199 225 1215
rect 159 1165 175 1199
rect 209 1165 225 1199
rect -15 1127 15 1149
rect 81 1127 111 1153
rect 159 1149 225 1165
rect 351 1199 417 1215
rect 351 1165 367 1199
rect 401 1165 417 1199
rect 177 1127 207 1149
rect 273 1127 303 1153
rect 351 1149 417 1165
rect 543 1199 609 1215
rect 543 1165 559 1199
rect 593 1165 609 1199
rect 369 1127 399 1149
rect 465 1127 495 1153
rect 543 1149 609 1165
rect 735 1199 801 1215
rect 735 1165 751 1199
rect 785 1165 801 1199
rect 561 1127 591 1149
rect 657 1127 687 1153
rect 735 1149 801 1165
rect 927 1199 993 1215
rect 927 1165 943 1199
rect 977 1165 993 1199
rect 753 1127 783 1149
rect 849 1127 879 1153
rect 927 1149 993 1165
rect 1119 1199 1185 1215
rect 1119 1165 1135 1199
rect 1169 1165 1185 1199
rect 945 1127 975 1149
rect 1041 1127 1071 1153
rect 1119 1149 1185 1165
rect 1137 1127 1167 1149
rect -1167 701 -1137 727
rect -1071 705 -1041 727
rect -1089 689 -1023 705
rect -975 701 -945 727
rect -879 705 -849 727
rect -1089 655 -1073 689
rect -1039 655 -1023 689
rect -1089 639 -1023 655
rect -897 689 -831 705
rect -783 701 -753 727
rect -687 705 -657 727
rect -897 655 -881 689
rect -847 655 -831 689
rect -897 639 -831 655
rect -705 689 -639 705
rect -591 701 -561 727
rect -495 705 -465 727
rect -705 655 -689 689
rect -655 655 -639 689
rect -705 639 -639 655
rect -513 689 -447 705
rect -399 701 -369 727
rect -303 705 -273 727
rect -513 655 -497 689
rect -463 655 -447 689
rect -513 639 -447 655
rect -321 689 -255 705
rect -207 701 -177 727
rect -111 705 -81 727
rect -321 655 -305 689
rect -271 655 -255 689
rect -321 639 -255 655
rect -129 689 -63 705
rect -15 701 15 727
rect 81 705 111 727
rect -129 655 -113 689
rect -79 655 -63 689
rect -129 639 -63 655
rect 63 689 129 705
rect 177 701 207 727
rect 273 705 303 727
rect 63 655 79 689
rect 113 655 129 689
rect 63 639 129 655
rect 255 689 321 705
rect 369 701 399 727
rect 465 705 495 727
rect 255 655 271 689
rect 305 655 321 689
rect 255 639 321 655
rect 447 689 513 705
rect 561 701 591 727
rect 657 705 687 727
rect 447 655 463 689
rect 497 655 513 689
rect 447 639 513 655
rect 639 689 705 705
rect 753 701 783 727
rect 849 705 879 727
rect 639 655 655 689
rect 689 655 705 689
rect 639 639 705 655
rect 831 689 897 705
rect 945 701 975 727
rect 1041 705 1071 727
rect 831 655 847 689
rect 881 655 897 689
rect 831 639 897 655
rect 1023 689 1089 705
rect 1137 701 1167 727
rect 1023 655 1039 689
rect 1073 655 1089 689
rect 1023 639 1089 655
rect -1089 581 -1023 597
rect -1089 547 -1073 581
rect -1039 547 -1023 581
rect -1167 509 -1137 535
rect -1089 531 -1023 547
rect -897 581 -831 597
rect -897 547 -881 581
rect -847 547 -831 581
rect -1071 509 -1041 531
rect -975 509 -945 535
rect -897 531 -831 547
rect -705 581 -639 597
rect -705 547 -689 581
rect -655 547 -639 581
rect -879 509 -849 531
rect -783 509 -753 535
rect -705 531 -639 547
rect -513 581 -447 597
rect -513 547 -497 581
rect -463 547 -447 581
rect -687 509 -657 531
rect -591 509 -561 535
rect -513 531 -447 547
rect -321 581 -255 597
rect -321 547 -305 581
rect -271 547 -255 581
rect -495 509 -465 531
rect -399 509 -369 535
rect -321 531 -255 547
rect -129 581 -63 597
rect -129 547 -113 581
rect -79 547 -63 581
rect -303 509 -273 531
rect -207 509 -177 535
rect -129 531 -63 547
rect 63 581 129 597
rect 63 547 79 581
rect 113 547 129 581
rect -111 509 -81 531
rect -15 509 15 535
rect 63 531 129 547
rect 255 581 321 597
rect 255 547 271 581
rect 305 547 321 581
rect 81 509 111 531
rect 177 509 207 535
rect 255 531 321 547
rect 447 581 513 597
rect 447 547 463 581
rect 497 547 513 581
rect 273 509 303 531
rect 369 509 399 535
rect 447 531 513 547
rect 639 581 705 597
rect 639 547 655 581
rect 689 547 705 581
rect 465 509 495 531
rect 561 509 591 535
rect 639 531 705 547
rect 831 581 897 597
rect 831 547 847 581
rect 881 547 897 581
rect 657 509 687 531
rect 753 509 783 535
rect 831 531 897 547
rect 1023 581 1089 597
rect 1023 547 1039 581
rect 1073 547 1089 581
rect 849 509 879 531
rect 945 509 975 535
rect 1023 531 1089 547
rect 1041 509 1071 531
rect 1137 509 1167 535
rect -1167 87 -1137 109
rect -1185 71 -1119 87
rect -1071 83 -1041 109
rect -975 87 -945 109
rect -1185 37 -1169 71
rect -1135 37 -1119 71
rect -1185 21 -1119 37
rect -993 71 -927 87
rect -879 83 -849 109
rect -783 87 -753 109
rect -993 37 -977 71
rect -943 37 -927 71
rect -993 21 -927 37
rect -801 71 -735 87
rect -687 83 -657 109
rect -591 87 -561 109
rect -801 37 -785 71
rect -751 37 -735 71
rect -801 21 -735 37
rect -609 71 -543 87
rect -495 83 -465 109
rect -399 87 -369 109
rect -609 37 -593 71
rect -559 37 -543 71
rect -609 21 -543 37
rect -417 71 -351 87
rect -303 83 -273 109
rect -207 87 -177 109
rect -417 37 -401 71
rect -367 37 -351 71
rect -417 21 -351 37
rect -225 71 -159 87
rect -111 83 -81 109
rect -15 87 15 109
rect -225 37 -209 71
rect -175 37 -159 71
rect -225 21 -159 37
rect -33 71 33 87
rect 81 83 111 109
rect 177 87 207 109
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 159 71 225 87
rect 273 83 303 109
rect 369 87 399 109
rect 159 37 175 71
rect 209 37 225 71
rect 159 21 225 37
rect 351 71 417 87
rect 465 83 495 109
rect 561 87 591 109
rect 351 37 367 71
rect 401 37 417 71
rect 351 21 417 37
rect 543 71 609 87
rect 657 83 687 109
rect 753 87 783 109
rect 543 37 559 71
rect 593 37 609 71
rect 543 21 609 37
rect 735 71 801 87
rect 849 83 879 109
rect 945 87 975 109
rect 735 37 751 71
rect 785 37 801 71
rect 735 21 801 37
rect 927 71 993 87
rect 1041 83 1071 109
rect 1137 87 1167 109
rect 927 37 943 71
rect 977 37 993 71
rect 927 21 993 37
rect 1119 71 1185 87
rect 1119 37 1135 71
rect 1169 37 1185 71
rect 1119 21 1185 37
rect -1185 -37 -1119 -21
rect -1185 -71 -1169 -37
rect -1135 -71 -1119 -37
rect -1185 -87 -1119 -71
rect -993 -37 -927 -21
rect -993 -71 -977 -37
rect -943 -71 -927 -37
rect -1167 -109 -1137 -87
rect -1071 -109 -1041 -83
rect -993 -87 -927 -71
rect -801 -37 -735 -21
rect -801 -71 -785 -37
rect -751 -71 -735 -37
rect -975 -109 -945 -87
rect -879 -109 -849 -83
rect -801 -87 -735 -71
rect -609 -37 -543 -21
rect -609 -71 -593 -37
rect -559 -71 -543 -37
rect -783 -109 -753 -87
rect -687 -109 -657 -83
rect -609 -87 -543 -71
rect -417 -37 -351 -21
rect -417 -71 -401 -37
rect -367 -71 -351 -37
rect -591 -109 -561 -87
rect -495 -109 -465 -83
rect -417 -87 -351 -71
rect -225 -37 -159 -21
rect -225 -71 -209 -37
rect -175 -71 -159 -37
rect -399 -109 -369 -87
rect -303 -109 -273 -83
rect -225 -87 -159 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -207 -109 -177 -87
rect -111 -109 -81 -83
rect -33 -87 33 -71
rect 159 -37 225 -21
rect 159 -71 175 -37
rect 209 -71 225 -37
rect -15 -109 15 -87
rect 81 -109 111 -83
rect 159 -87 225 -71
rect 351 -37 417 -21
rect 351 -71 367 -37
rect 401 -71 417 -37
rect 177 -109 207 -87
rect 273 -109 303 -83
rect 351 -87 417 -71
rect 543 -37 609 -21
rect 543 -71 559 -37
rect 593 -71 609 -37
rect 369 -109 399 -87
rect 465 -109 495 -83
rect 543 -87 609 -71
rect 735 -37 801 -21
rect 735 -71 751 -37
rect 785 -71 801 -37
rect 561 -109 591 -87
rect 657 -109 687 -83
rect 735 -87 801 -71
rect 927 -37 993 -21
rect 927 -71 943 -37
rect 977 -71 993 -37
rect 753 -109 783 -87
rect 849 -109 879 -83
rect 927 -87 993 -71
rect 1119 -37 1185 -21
rect 1119 -71 1135 -37
rect 1169 -71 1185 -37
rect 945 -109 975 -87
rect 1041 -109 1071 -83
rect 1119 -87 1185 -71
rect 1137 -109 1167 -87
rect -1167 -535 -1137 -509
rect -1071 -531 -1041 -509
rect -1089 -547 -1023 -531
rect -975 -535 -945 -509
rect -879 -531 -849 -509
rect -1089 -581 -1073 -547
rect -1039 -581 -1023 -547
rect -1089 -597 -1023 -581
rect -897 -547 -831 -531
rect -783 -535 -753 -509
rect -687 -531 -657 -509
rect -897 -581 -881 -547
rect -847 -581 -831 -547
rect -897 -597 -831 -581
rect -705 -547 -639 -531
rect -591 -535 -561 -509
rect -495 -531 -465 -509
rect -705 -581 -689 -547
rect -655 -581 -639 -547
rect -705 -597 -639 -581
rect -513 -547 -447 -531
rect -399 -535 -369 -509
rect -303 -531 -273 -509
rect -513 -581 -497 -547
rect -463 -581 -447 -547
rect -513 -597 -447 -581
rect -321 -547 -255 -531
rect -207 -535 -177 -509
rect -111 -531 -81 -509
rect -321 -581 -305 -547
rect -271 -581 -255 -547
rect -321 -597 -255 -581
rect -129 -547 -63 -531
rect -15 -535 15 -509
rect 81 -531 111 -509
rect -129 -581 -113 -547
rect -79 -581 -63 -547
rect -129 -597 -63 -581
rect 63 -547 129 -531
rect 177 -535 207 -509
rect 273 -531 303 -509
rect 63 -581 79 -547
rect 113 -581 129 -547
rect 63 -597 129 -581
rect 255 -547 321 -531
rect 369 -535 399 -509
rect 465 -531 495 -509
rect 255 -581 271 -547
rect 305 -581 321 -547
rect 255 -597 321 -581
rect 447 -547 513 -531
rect 561 -535 591 -509
rect 657 -531 687 -509
rect 447 -581 463 -547
rect 497 -581 513 -547
rect 447 -597 513 -581
rect 639 -547 705 -531
rect 753 -535 783 -509
rect 849 -531 879 -509
rect 639 -581 655 -547
rect 689 -581 705 -547
rect 639 -597 705 -581
rect 831 -547 897 -531
rect 945 -535 975 -509
rect 1041 -531 1071 -509
rect 831 -581 847 -547
rect 881 -581 897 -547
rect 831 -597 897 -581
rect 1023 -547 1089 -531
rect 1137 -535 1167 -509
rect 1023 -581 1039 -547
rect 1073 -581 1089 -547
rect 1023 -597 1089 -581
rect -1089 -655 -1023 -639
rect -1089 -689 -1073 -655
rect -1039 -689 -1023 -655
rect -1167 -727 -1137 -701
rect -1089 -705 -1023 -689
rect -897 -655 -831 -639
rect -897 -689 -881 -655
rect -847 -689 -831 -655
rect -1071 -727 -1041 -705
rect -975 -727 -945 -701
rect -897 -705 -831 -689
rect -705 -655 -639 -639
rect -705 -689 -689 -655
rect -655 -689 -639 -655
rect -879 -727 -849 -705
rect -783 -727 -753 -701
rect -705 -705 -639 -689
rect -513 -655 -447 -639
rect -513 -689 -497 -655
rect -463 -689 -447 -655
rect -687 -727 -657 -705
rect -591 -727 -561 -701
rect -513 -705 -447 -689
rect -321 -655 -255 -639
rect -321 -689 -305 -655
rect -271 -689 -255 -655
rect -495 -727 -465 -705
rect -399 -727 -369 -701
rect -321 -705 -255 -689
rect -129 -655 -63 -639
rect -129 -689 -113 -655
rect -79 -689 -63 -655
rect -303 -727 -273 -705
rect -207 -727 -177 -701
rect -129 -705 -63 -689
rect 63 -655 129 -639
rect 63 -689 79 -655
rect 113 -689 129 -655
rect -111 -727 -81 -705
rect -15 -727 15 -701
rect 63 -705 129 -689
rect 255 -655 321 -639
rect 255 -689 271 -655
rect 305 -689 321 -655
rect 81 -727 111 -705
rect 177 -727 207 -701
rect 255 -705 321 -689
rect 447 -655 513 -639
rect 447 -689 463 -655
rect 497 -689 513 -655
rect 273 -727 303 -705
rect 369 -727 399 -701
rect 447 -705 513 -689
rect 639 -655 705 -639
rect 639 -689 655 -655
rect 689 -689 705 -655
rect 465 -727 495 -705
rect 561 -727 591 -701
rect 639 -705 705 -689
rect 831 -655 897 -639
rect 831 -689 847 -655
rect 881 -689 897 -655
rect 657 -727 687 -705
rect 753 -727 783 -701
rect 831 -705 897 -689
rect 1023 -655 1089 -639
rect 1023 -689 1039 -655
rect 1073 -689 1089 -655
rect 849 -727 879 -705
rect 945 -727 975 -701
rect 1023 -705 1089 -689
rect 1041 -727 1071 -705
rect 1137 -727 1167 -701
rect -1167 -1149 -1137 -1127
rect -1185 -1165 -1119 -1149
rect -1071 -1153 -1041 -1127
rect -975 -1149 -945 -1127
rect -1185 -1199 -1169 -1165
rect -1135 -1199 -1119 -1165
rect -1185 -1215 -1119 -1199
rect -993 -1165 -927 -1149
rect -879 -1153 -849 -1127
rect -783 -1149 -753 -1127
rect -993 -1199 -977 -1165
rect -943 -1199 -927 -1165
rect -993 -1215 -927 -1199
rect -801 -1165 -735 -1149
rect -687 -1153 -657 -1127
rect -591 -1149 -561 -1127
rect -801 -1199 -785 -1165
rect -751 -1199 -735 -1165
rect -801 -1215 -735 -1199
rect -609 -1165 -543 -1149
rect -495 -1153 -465 -1127
rect -399 -1149 -369 -1127
rect -609 -1199 -593 -1165
rect -559 -1199 -543 -1165
rect -609 -1215 -543 -1199
rect -417 -1165 -351 -1149
rect -303 -1153 -273 -1127
rect -207 -1149 -177 -1127
rect -417 -1199 -401 -1165
rect -367 -1199 -351 -1165
rect -417 -1215 -351 -1199
rect -225 -1165 -159 -1149
rect -111 -1153 -81 -1127
rect -15 -1149 15 -1127
rect -225 -1199 -209 -1165
rect -175 -1199 -159 -1165
rect -225 -1215 -159 -1199
rect -33 -1165 33 -1149
rect 81 -1153 111 -1127
rect 177 -1149 207 -1127
rect -33 -1199 -17 -1165
rect 17 -1199 33 -1165
rect -33 -1215 33 -1199
rect 159 -1165 225 -1149
rect 273 -1153 303 -1127
rect 369 -1149 399 -1127
rect 159 -1199 175 -1165
rect 209 -1199 225 -1165
rect 159 -1215 225 -1199
rect 351 -1165 417 -1149
rect 465 -1153 495 -1127
rect 561 -1149 591 -1127
rect 351 -1199 367 -1165
rect 401 -1199 417 -1165
rect 351 -1215 417 -1199
rect 543 -1165 609 -1149
rect 657 -1153 687 -1127
rect 753 -1149 783 -1127
rect 543 -1199 559 -1165
rect 593 -1199 609 -1165
rect 543 -1215 609 -1199
rect 735 -1165 801 -1149
rect 849 -1153 879 -1127
rect 945 -1149 975 -1127
rect 735 -1199 751 -1165
rect 785 -1199 801 -1165
rect 735 -1215 801 -1199
rect 927 -1165 993 -1149
rect 1041 -1153 1071 -1127
rect 1137 -1149 1167 -1127
rect 927 -1199 943 -1165
rect 977 -1199 993 -1165
rect 927 -1215 993 -1199
rect 1119 -1165 1185 -1149
rect 1119 -1199 1135 -1165
rect 1169 -1199 1185 -1165
rect 1119 -1215 1185 -1199
<< polycont >>
rect -1169 1165 -1135 1199
rect -977 1165 -943 1199
rect -785 1165 -751 1199
rect -593 1165 -559 1199
rect -401 1165 -367 1199
rect -209 1165 -175 1199
rect -17 1165 17 1199
rect 175 1165 209 1199
rect 367 1165 401 1199
rect 559 1165 593 1199
rect 751 1165 785 1199
rect 943 1165 977 1199
rect 1135 1165 1169 1199
rect -1073 655 -1039 689
rect -881 655 -847 689
rect -689 655 -655 689
rect -497 655 -463 689
rect -305 655 -271 689
rect -113 655 -79 689
rect 79 655 113 689
rect 271 655 305 689
rect 463 655 497 689
rect 655 655 689 689
rect 847 655 881 689
rect 1039 655 1073 689
rect -1073 547 -1039 581
rect -881 547 -847 581
rect -689 547 -655 581
rect -497 547 -463 581
rect -305 547 -271 581
rect -113 547 -79 581
rect 79 547 113 581
rect 271 547 305 581
rect 463 547 497 581
rect 655 547 689 581
rect 847 547 881 581
rect 1039 547 1073 581
rect -1169 37 -1135 71
rect -977 37 -943 71
rect -785 37 -751 71
rect -593 37 -559 71
rect -401 37 -367 71
rect -209 37 -175 71
rect -17 37 17 71
rect 175 37 209 71
rect 367 37 401 71
rect 559 37 593 71
rect 751 37 785 71
rect 943 37 977 71
rect 1135 37 1169 71
rect -1169 -71 -1135 -37
rect -977 -71 -943 -37
rect -785 -71 -751 -37
rect -593 -71 -559 -37
rect -401 -71 -367 -37
rect -209 -71 -175 -37
rect -17 -71 17 -37
rect 175 -71 209 -37
rect 367 -71 401 -37
rect 559 -71 593 -37
rect 751 -71 785 -37
rect 943 -71 977 -37
rect 1135 -71 1169 -37
rect -1073 -581 -1039 -547
rect -881 -581 -847 -547
rect -689 -581 -655 -547
rect -497 -581 -463 -547
rect -305 -581 -271 -547
rect -113 -581 -79 -547
rect 79 -581 113 -547
rect 271 -581 305 -547
rect 463 -581 497 -547
rect 655 -581 689 -547
rect 847 -581 881 -547
rect 1039 -581 1073 -547
rect -1073 -689 -1039 -655
rect -881 -689 -847 -655
rect -689 -689 -655 -655
rect -497 -689 -463 -655
rect -305 -689 -271 -655
rect -113 -689 -79 -655
rect 79 -689 113 -655
rect 271 -689 305 -655
rect 463 -689 497 -655
rect 655 -689 689 -655
rect 847 -689 881 -655
rect 1039 -689 1073 -655
rect -1169 -1199 -1135 -1165
rect -977 -1199 -943 -1165
rect -785 -1199 -751 -1165
rect -593 -1199 -559 -1165
rect -401 -1199 -367 -1165
rect -209 -1199 -175 -1165
rect -17 -1199 17 -1165
rect 175 -1199 209 -1165
rect 367 -1199 401 -1165
rect 559 -1199 593 -1165
rect 751 -1199 785 -1165
rect 943 -1199 977 -1165
rect 1135 -1199 1169 -1165
<< locali >>
rect -1331 1267 -1235 1301
rect 1235 1267 1331 1301
rect -1331 1205 -1297 1267
rect 1297 1205 1331 1267
rect -1185 1165 -1169 1199
rect -1135 1165 -1119 1199
rect -993 1165 -977 1199
rect -943 1165 -927 1199
rect -801 1165 -785 1199
rect -751 1165 -735 1199
rect -609 1165 -593 1199
rect -559 1165 -543 1199
rect -417 1165 -401 1199
rect -367 1165 -351 1199
rect -225 1165 -209 1199
rect -175 1165 -159 1199
rect -33 1165 -17 1199
rect 17 1165 33 1199
rect 159 1165 175 1199
rect 209 1165 225 1199
rect 351 1165 367 1199
rect 401 1165 417 1199
rect 543 1165 559 1199
rect 593 1165 609 1199
rect 735 1165 751 1199
rect 785 1165 801 1199
rect 927 1165 943 1199
rect 977 1165 993 1199
rect 1119 1165 1135 1199
rect 1169 1165 1185 1199
rect -1217 1115 -1183 1131
rect -1217 723 -1183 739
rect -1121 1115 -1087 1131
rect -1121 723 -1087 739
rect -1025 1115 -991 1131
rect -1025 723 -991 739
rect -929 1115 -895 1131
rect -929 723 -895 739
rect -833 1115 -799 1131
rect -833 723 -799 739
rect -737 1115 -703 1131
rect -737 723 -703 739
rect -641 1115 -607 1131
rect -641 723 -607 739
rect -545 1115 -511 1131
rect -545 723 -511 739
rect -449 1115 -415 1131
rect -449 723 -415 739
rect -353 1115 -319 1131
rect -353 723 -319 739
rect -257 1115 -223 1131
rect -257 723 -223 739
rect -161 1115 -127 1131
rect -161 723 -127 739
rect -65 1115 -31 1131
rect -65 723 -31 739
rect 31 1115 65 1131
rect 31 723 65 739
rect 127 1115 161 1131
rect 127 723 161 739
rect 223 1115 257 1131
rect 223 723 257 739
rect 319 1115 353 1131
rect 319 723 353 739
rect 415 1115 449 1131
rect 415 723 449 739
rect 511 1115 545 1131
rect 511 723 545 739
rect 607 1115 641 1131
rect 607 723 641 739
rect 703 1115 737 1131
rect 703 723 737 739
rect 799 1115 833 1131
rect 799 723 833 739
rect 895 1115 929 1131
rect 895 723 929 739
rect 991 1115 1025 1131
rect 991 723 1025 739
rect 1087 1115 1121 1131
rect 1087 723 1121 739
rect 1183 1115 1217 1131
rect 1183 723 1217 739
rect -1089 655 -1073 689
rect -1039 655 -1023 689
rect -897 655 -881 689
rect -847 655 -831 689
rect -705 655 -689 689
rect -655 655 -639 689
rect -513 655 -497 689
rect -463 655 -447 689
rect -321 655 -305 689
rect -271 655 -255 689
rect -129 655 -113 689
rect -79 655 -63 689
rect 63 655 79 689
rect 113 655 129 689
rect 255 655 271 689
rect 305 655 321 689
rect 447 655 463 689
rect 497 655 513 689
rect 639 655 655 689
rect 689 655 705 689
rect 831 655 847 689
rect 881 655 897 689
rect 1023 655 1039 689
rect 1073 655 1089 689
rect -1089 547 -1073 581
rect -1039 547 -1023 581
rect -897 547 -881 581
rect -847 547 -831 581
rect -705 547 -689 581
rect -655 547 -639 581
rect -513 547 -497 581
rect -463 547 -447 581
rect -321 547 -305 581
rect -271 547 -255 581
rect -129 547 -113 581
rect -79 547 -63 581
rect 63 547 79 581
rect 113 547 129 581
rect 255 547 271 581
rect 305 547 321 581
rect 447 547 463 581
rect 497 547 513 581
rect 639 547 655 581
rect 689 547 705 581
rect 831 547 847 581
rect 881 547 897 581
rect 1023 547 1039 581
rect 1073 547 1089 581
rect -1217 497 -1183 513
rect -1217 105 -1183 121
rect -1121 497 -1087 513
rect -1121 105 -1087 121
rect -1025 497 -991 513
rect -1025 105 -991 121
rect -929 497 -895 513
rect -929 105 -895 121
rect -833 497 -799 513
rect -833 105 -799 121
rect -737 497 -703 513
rect -737 105 -703 121
rect -641 497 -607 513
rect -641 105 -607 121
rect -545 497 -511 513
rect -545 105 -511 121
rect -449 497 -415 513
rect -449 105 -415 121
rect -353 497 -319 513
rect -353 105 -319 121
rect -257 497 -223 513
rect -257 105 -223 121
rect -161 497 -127 513
rect -161 105 -127 121
rect -65 497 -31 513
rect -65 105 -31 121
rect 31 497 65 513
rect 31 105 65 121
rect 127 497 161 513
rect 127 105 161 121
rect 223 497 257 513
rect 223 105 257 121
rect 319 497 353 513
rect 319 105 353 121
rect 415 497 449 513
rect 415 105 449 121
rect 511 497 545 513
rect 511 105 545 121
rect 607 497 641 513
rect 607 105 641 121
rect 703 497 737 513
rect 703 105 737 121
rect 799 497 833 513
rect 799 105 833 121
rect 895 497 929 513
rect 895 105 929 121
rect 991 497 1025 513
rect 991 105 1025 121
rect 1087 497 1121 513
rect 1087 105 1121 121
rect 1183 497 1217 513
rect 1183 105 1217 121
rect -1185 37 -1169 71
rect -1135 37 -1119 71
rect -993 37 -977 71
rect -943 37 -927 71
rect -801 37 -785 71
rect -751 37 -735 71
rect -609 37 -593 71
rect -559 37 -543 71
rect -417 37 -401 71
rect -367 37 -351 71
rect -225 37 -209 71
rect -175 37 -159 71
rect -33 37 -17 71
rect 17 37 33 71
rect 159 37 175 71
rect 209 37 225 71
rect 351 37 367 71
rect 401 37 417 71
rect 543 37 559 71
rect 593 37 609 71
rect 735 37 751 71
rect 785 37 801 71
rect 927 37 943 71
rect 977 37 993 71
rect 1119 37 1135 71
rect 1169 37 1185 71
rect -1185 -71 -1169 -37
rect -1135 -71 -1119 -37
rect -993 -71 -977 -37
rect -943 -71 -927 -37
rect -801 -71 -785 -37
rect -751 -71 -735 -37
rect -609 -71 -593 -37
rect -559 -71 -543 -37
rect -417 -71 -401 -37
rect -367 -71 -351 -37
rect -225 -71 -209 -37
rect -175 -71 -159 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 159 -71 175 -37
rect 209 -71 225 -37
rect 351 -71 367 -37
rect 401 -71 417 -37
rect 543 -71 559 -37
rect 593 -71 609 -37
rect 735 -71 751 -37
rect 785 -71 801 -37
rect 927 -71 943 -37
rect 977 -71 993 -37
rect 1119 -71 1135 -37
rect 1169 -71 1185 -37
rect -1217 -121 -1183 -105
rect -1217 -513 -1183 -497
rect -1121 -121 -1087 -105
rect -1121 -513 -1087 -497
rect -1025 -121 -991 -105
rect -1025 -513 -991 -497
rect -929 -121 -895 -105
rect -929 -513 -895 -497
rect -833 -121 -799 -105
rect -833 -513 -799 -497
rect -737 -121 -703 -105
rect -737 -513 -703 -497
rect -641 -121 -607 -105
rect -641 -513 -607 -497
rect -545 -121 -511 -105
rect -545 -513 -511 -497
rect -449 -121 -415 -105
rect -449 -513 -415 -497
rect -353 -121 -319 -105
rect -353 -513 -319 -497
rect -257 -121 -223 -105
rect -257 -513 -223 -497
rect -161 -121 -127 -105
rect -161 -513 -127 -497
rect -65 -121 -31 -105
rect -65 -513 -31 -497
rect 31 -121 65 -105
rect 31 -513 65 -497
rect 127 -121 161 -105
rect 127 -513 161 -497
rect 223 -121 257 -105
rect 223 -513 257 -497
rect 319 -121 353 -105
rect 319 -513 353 -497
rect 415 -121 449 -105
rect 415 -513 449 -497
rect 511 -121 545 -105
rect 511 -513 545 -497
rect 607 -121 641 -105
rect 607 -513 641 -497
rect 703 -121 737 -105
rect 703 -513 737 -497
rect 799 -121 833 -105
rect 799 -513 833 -497
rect 895 -121 929 -105
rect 895 -513 929 -497
rect 991 -121 1025 -105
rect 991 -513 1025 -497
rect 1087 -121 1121 -105
rect 1087 -513 1121 -497
rect 1183 -121 1217 -105
rect 1183 -513 1217 -497
rect -1089 -581 -1073 -547
rect -1039 -581 -1023 -547
rect -897 -581 -881 -547
rect -847 -581 -831 -547
rect -705 -581 -689 -547
rect -655 -581 -639 -547
rect -513 -581 -497 -547
rect -463 -581 -447 -547
rect -321 -581 -305 -547
rect -271 -581 -255 -547
rect -129 -581 -113 -547
rect -79 -581 -63 -547
rect 63 -581 79 -547
rect 113 -581 129 -547
rect 255 -581 271 -547
rect 305 -581 321 -547
rect 447 -581 463 -547
rect 497 -581 513 -547
rect 639 -581 655 -547
rect 689 -581 705 -547
rect 831 -581 847 -547
rect 881 -581 897 -547
rect 1023 -581 1039 -547
rect 1073 -581 1089 -547
rect -1089 -689 -1073 -655
rect -1039 -689 -1023 -655
rect -897 -689 -881 -655
rect -847 -689 -831 -655
rect -705 -689 -689 -655
rect -655 -689 -639 -655
rect -513 -689 -497 -655
rect -463 -689 -447 -655
rect -321 -689 -305 -655
rect -271 -689 -255 -655
rect -129 -689 -113 -655
rect -79 -689 -63 -655
rect 63 -689 79 -655
rect 113 -689 129 -655
rect 255 -689 271 -655
rect 305 -689 321 -655
rect 447 -689 463 -655
rect 497 -689 513 -655
rect 639 -689 655 -655
rect 689 -689 705 -655
rect 831 -689 847 -655
rect 881 -689 897 -655
rect 1023 -689 1039 -655
rect 1073 -689 1089 -655
rect -1217 -739 -1183 -723
rect -1217 -1131 -1183 -1115
rect -1121 -739 -1087 -723
rect -1121 -1131 -1087 -1115
rect -1025 -739 -991 -723
rect -1025 -1131 -991 -1115
rect -929 -739 -895 -723
rect -929 -1131 -895 -1115
rect -833 -739 -799 -723
rect -833 -1131 -799 -1115
rect -737 -739 -703 -723
rect -737 -1131 -703 -1115
rect -641 -739 -607 -723
rect -641 -1131 -607 -1115
rect -545 -739 -511 -723
rect -545 -1131 -511 -1115
rect -449 -739 -415 -723
rect -449 -1131 -415 -1115
rect -353 -739 -319 -723
rect -353 -1131 -319 -1115
rect -257 -739 -223 -723
rect -257 -1131 -223 -1115
rect -161 -739 -127 -723
rect -161 -1131 -127 -1115
rect -65 -739 -31 -723
rect -65 -1131 -31 -1115
rect 31 -739 65 -723
rect 31 -1131 65 -1115
rect 127 -739 161 -723
rect 127 -1131 161 -1115
rect 223 -739 257 -723
rect 223 -1131 257 -1115
rect 319 -739 353 -723
rect 319 -1131 353 -1115
rect 415 -739 449 -723
rect 415 -1131 449 -1115
rect 511 -739 545 -723
rect 511 -1131 545 -1115
rect 607 -739 641 -723
rect 607 -1131 641 -1115
rect 703 -739 737 -723
rect 703 -1131 737 -1115
rect 799 -739 833 -723
rect 799 -1131 833 -1115
rect 895 -739 929 -723
rect 895 -1131 929 -1115
rect 991 -739 1025 -723
rect 991 -1131 1025 -1115
rect 1087 -739 1121 -723
rect 1087 -1131 1121 -1115
rect 1183 -739 1217 -723
rect 1183 -1131 1217 -1115
rect -1185 -1199 -1169 -1165
rect -1135 -1199 -1119 -1165
rect -993 -1199 -977 -1165
rect -943 -1199 -927 -1165
rect -801 -1199 -785 -1165
rect -751 -1199 -735 -1165
rect -609 -1199 -593 -1165
rect -559 -1199 -543 -1165
rect -417 -1199 -401 -1165
rect -367 -1199 -351 -1165
rect -225 -1199 -209 -1165
rect -175 -1199 -159 -1165
rect -33 -1199 -17 -1165
rect 17 -1199 33 -1165
rect 159 -1199 175 -1165
rect 209 -1199 225 -1165
rect 351 -1199 367 -1165
rect 401 -1199 417 -1165
rect 543 -1199 559 -1165
rect 593 -1199 609 -1165
rect 735 -1199 751 -1165
rect 785 -1199 801 -1165
rect 927 -1199 943 -1165
rect 977 -1199 993 -1165
rect 1119 -1199 1135 -1165
rect 1169 -1199 1185 -1165
rect -1331 -1267 -1297 -1205
rect 1297 -1267 1331 -1205
rect -1331 -1301 -1235 -1267
rect 1235 -1301 1331 -1267
<< viali >>
rect -1169 1165 -1135 1199
rect -977 1165 -943 1199
rect -785 1165 -751 1199
rect -593 1165 -559 1199
rect -401 1165 -367 1199
rect -209 1165 -175 1199
rect -17 1165 17 1199
rect 175 1165 209 1199
rect 367 1165 401 1199
rect 559 1165 593 1199
rect 751 1165 785 1199
rect 943 1165 977 1199
rect 1135 1165 1169 1199
rect -1217 739 -1183 1115
rect -1121 739 -1087 1115
rect -1025 739 -991 1115
rect -929 739 -895 1115
rect -833 739 -799 1115
rect -737 739 -703 1115
rect -641 739 -607 1115
rect -545 739 -511 1115
rect -449 739 -415 1115
rect -353 739 -319 1115
rect -257 739 -223 1115
rect -161 739 -127 1115
rect -65 739 -31 1115
rect 31 739 65 1115
rect 127 739 161 1115
rect 223 739 257 1115
rect 319 739 353 1115
rect 415 739 449 1115
rect 511 739 545 1115
rect 607 739 641 1115
rect 703 739 737 1115
rect 799 739 833 1115
rect 895 739 929 1115
rect 991 739 1025 1115
rect 1087 739 1121 1115
rect 1183 739 1217 1115
rect -1073 655 -1039 689
rect -881 655 -847 689
rect -689 655 -655 689
rect -497 655 -463 689
rect -305 655 -271 689
rect -113 655 -79 689
rect 79 655 113 689
rect 271 655 305 689
rect 463 655 497 689
rect 655 655 689 689
rect 847 655 881 689
rect 1039 655 1073 689
rect -1073 547 -1039 581
rect -881 547 -847 581
rect -689 547 -655 581
rect -497 547 -463 581
rect -305 547 -271 581
rect -113 547 -79 581
rect 79 547 113 581
rect 271 547 305 581
rect 463 547 497 581
rect 655 547 689 581
rect 847 547 881 581
rect 1039 547 1073 581
rect -1217 121 -1183 497
rect -1121 121 -1087 497
rect -1025 121 -991 497
rect -929 121 -895 497
rect -833 121 -799 497
rect -737 121 -703 497
rect -641 121 -607 497
rect -545 121 -511 497
rect -449 121 -415 497
rect -353 121 -319 497
rect -257 121 -223 497
rect -161 121 -127 497
rect -65 121 -31 497
rect 31 121 65 497
rect 127 121 161 497
rect 223 121 257 497
rect 319 121 353 497
rect 415 121 449 497
rect 511 121 545 497
rect 607 121 641 497
rect 703 121 737 497
rect 799 121 833 497
rect 895 121 929 497
rect 991 121 1025 497
rect 1087 121 1121 497
rect 1183 121 1217 497
rect -1169 37 -1135 71
rect -977 37 -943 71
rect -785 37 -751 71
rect -593 37 -559 71
rect -401 37 -367 71
rect -209 37 -175 71
rect -17 37 17 71
rect 175 37 209 71
rect 367 37 401 71
rect 559 37 593 71
rect 751 37 785 71
rect 943 37 977 71
rect 1135 37 1169 71
rect -1169 -71 -1135 -37
rect -977 -71 -943 -37
rect -785 -71 -751 -37
rect -593 -71 -559 -37
rect -401 -71 -367 -37
rect -209 -71 -175 -37
rect -17 -71 17 -37
rect 175 -71 209 -37
rect 367 -71 401 -37
rect 559 -71 593 -37
rect 751 -71 785 -37
rect 943 -71 977 -37
rect 1135 -71 1169 -37
rect -1217 -497 -1183 -121
rect -1121 -497 -1087 -121
rect -1025 -497 -991 -121
rect -929 -497 -895 -121
rect -833 -497 -799 -121
rect -737 -497 -703 -121
rect -641 -497 -607 -121
rect -545 -497 -511 -121
rect -449 -497 -415 -121
rect -353 -497 -319 -121
rect -257 -497 -223 -121
rect -161 -497 -127 -121
rect -65 -497 -31 -121
rect 31 -497 65 -121
rect 127 -497 161 -121
rect 223 -497 257 -121
rect 319 -497 353 -121
rect 415 -497 449 -121
rect 511 -497 545 -121
rect 607 -497 641 -121
rect 703 -497 737 -121
rect 799 -497 833 -121
rect 895 -497 929 -121
rect 991 -497 1025 -121
rect 1087 -497 1121 -121
rect 1183 -497 1217 -121
rect -1073 -581 -1039 -547
rect -881 -581 -847 -547
rect -689 -581 -655 -547
rect -497 -581 -463 -547
rect -305 -581 -271 -547
rect -113 -581 -79 -547
rect 79 -581 113 -547
rect 271 -581 305 -547
rect 463 -581 497 -547
rect 655 -581 689 -547
rect 847 -581 881 -547
rect 1039 -581 1073 -547
rect -1073 -689 -1039 -655
rect -881 -689 -847 -655
rect -689 -689 -655 -655
rect -497 -689 -463 -655
rect -305 -689 -271 -655
rect -113 -689 -79 -655
rect 79 -689 113 -655
rect 271 -689 305 -655
rect 463 -689 497 -655
rect 655 -689 689 -655
rect 847 -689 881 -655
rect 1039 -689 1073 -655
rect -1217 -1115 -1183 -739
rect -1121 -1115 -1087 -739
rect -1025 -1115 -991 -739
rect -929 -1115 -895 -739
rect -833 -1115 -799 -739
rect -737 -1115 -703 -739
rect -641 -1115 -607 -739
rect -545 -1115 -511 -739
rect -449 -1115 -415 -739
rect -353 -1115 -319 -739
rect -257 -1115 -223 -739
rect -161 -1115 -127 -739
rect -65 -1115 -31 -739
rect 31 -1115 65 -739
rect 127 -1115 161 -739
rect 223 -1115 257 -739
rect 319 -1115 353 -739
rect 415 -1115 449 -739
rect 511 -1115 545 -739
rect 607 -1115 641 -739
rect 703 -1115 737 -739
rect 799 -1115 833 -739
rect 895 -1115 929 -739
rect 991 -1115 1025 -739
rect 1087 -1115 1121 -739
rect 1183 -1115 1217 -739
rect -1169 -1199 -1135 -1165
rect -977 -1199 -943 -1165
rect -785 -1199 -751 -1165
rect -593 -1199 -559 -1165
rect -401 -1199 -367 -1165
rect -209 -1199 -175 -1165
rect -17 -1199 17 -1165
rect 175 -1199 209 -1165
rect 367 -1199 401 -1165
rect 559 -1199 593 -1165
rect 751 -1199 785 -1165
rect 943 -1199 977 -1165
rect 1135 -1199 1169 -1165
<< metal1 >>
rect -1181 1199 -1123 1205
rect -1181 1165 -1169 1199
rect -1135 1165 -1123 1199
rect -1181 1159 -1123 1165
rect -989 1199 -931 1205
rect -989 1165 -977 1199
rect -943 1165 -931 1199
rect -989 1159 -931 1165
rect -797 1199 -739 1205
rect -797 1165 -785 1199
rect -751 1165 -739 1199
rect -797 1159 -739 1165
rect -605 1199 -547 1205
rect -605 1165 -593 1199
rect -559 1165 -547 1199
rect -605 1159 -547 1165
rect -413 1199 -355 1205
rect -413 1165 -401 1199
rect -367 1165 -355 1199
rect -413 1159 -355 1165
rect -221 1199 -163 1205
rect -221 1165 -209 1199
rect -175 1165 -163 1199
rect -221 1159 -163 1165
rect -29 1199 29 1205
rect -29 1165 -17 1199
rect 17 1165 29 1199
rect -29 1159 29 1165
rect 163 1199 221 1205
rect 163 1165 175 1199
rect 209 1165 221 1199
rect 163 1159 221 1165
rect 355 1199 413 1205
rect 355 1165 367 1199
rect 401 1165 413 1199
rect 355 1159 413 1165
rect 547 1199 605 1205
rect 547 1165 559 1199
rect 593 1165 605 1199
rect 547 1159 605 1165
rect 739 1199 797 1205
rect 739 1165 751 1199
rect 785 1165 797 1199
rect 739 1159 797 1165
rect 931 1199 989 1205
rect 931 1165 943 1199
rect 977 1165 989 1199
rect 931 1159 989 1165
rect 1123 1199 1181 1205
rect 1123 1165 1135 1199
rect 1169 1165 1181 1199
rect 1123 1159 1181 1165
rect -1223 1115 -1177 1127
rect -1223 739 -1217 1115
rect -1183 739 -1177 1115
rect -1223 727 -1177 739
rect -1127 1115 -1081 1127
rect -1127 739 -1121 1115
rect -1087 739 -1081 1115
rect -1127 727 -1081 739
rect -1031 1115 -985 1127
rect -1031 739 -1025 1115
rect -991 739 -985 1115
rect -1031 727 -985 739
rect -935 1115 -889 1127
rect -935 739 -929 1115
rect -895 739 -889 1115
rect -935 727 -889 739
rect -839 1115 -793 1127
rect -839 739 -833 1115
rect -799 739 -793 1115
rect -839 727 -793 739
rect -743 1115 -697 1127
rect -743 739 -737 1115
rect -703 739 -697 1115
rect -743 727 -697 739
rect -647 1115 -601 1127
rect -647 739 -641 1115
rect -607 739 -601 1115
rect -647 727 -601 739
rect -551 1115 -505 1127
rect -551 739 -545 1115
rect -511 739 -505 1115
rect -551 727 -505 739
rect -455 1115 -409 1127
rect -455 739 -449 1115
rect -415 739 -409 1115
rect -455 727 -409 739
rect -359 1115 -313 1127
rect -359 739 -353 1115
rect -319 739 -313 1115
rect -359 727 -313 739
rect -263 1115 -217 1127
rect -263 739 -257 1115
rect -223 739 -217 1115
rect -263 727 -217 739
rect -167 1115 -121 1127
rect -167 739 -161 1115
rect -127 739 -121 1115
rect -167 727 -121 739
rect -71 1115 -25 1127
rect -71 739 -65 1115
rect -31 739 -25 1115
rect -71 727 -25 739
rect 25 1115 71 1127
rect 25 739 31 1115
rect 65 739 71 1115
rect 25 727 71 739
rect 121 1115 167 1127
rect 121 739 127 1115
rect 161 739 167 1115
rect 121 727 167 739
rect 217 1115 263 1127
rect 217 739 223 1115
rect 257 739 263 1115
rect 217 727 263 739
rect 313 1115 359 1127
rect 313 739 319 1115
rect 353 739 359 1115
rect 313 727 359 739
rect 409 1115 455 1127
rect 409 739 415 1115
rect 449 739 455 1115
rect 409 727 455 739
rect 505 1115 551 1127
rect 505 739 511 1115
rect 545 739 551 1115
rect 505 727 551 739
rect 601 1115 647 1127
rect 601 739 607 1115
rect 641 739 647 1115
rect 601 727 647 739
rect 697 1115 743 1127
rect 697 739 703 1115
rect 737 739 743 1115
rect 697 727 743 739
rect 793 1115 839 1127
rect 793 739 799 1115
rect 833 739 839 1115
rect 793 727 839 739
rect 889 1115 935 1127
rect 889 739 895 1115
rect 929 739 935 1115
rect 889 727 935 739
rect 985 1115 1031 1127
rect 985 739 991 1115
rect 1025 739 1031 1115
rect 985 727 1031 739
rect 1081 1115 1127 1127
rect 1081 739 1087 1115
rect 1121 739 1127 1115
rect 1081 727 1127 739
rect 1177 1115 1223 1127
rect 1177 739 1183 1115
rect 1217 739 1223 1115
rect 1177 727 1223 739
rect -1085 689 -1027 695
rect -1085 655 -1073 689
rect -1039 655 -1027 689
rect -1085 649 -1027 655
rect -893 689 -835 695
rect -893 655 -881 689
rect -847 655 -835 689
rect -893 649 -835 655
rect -701 689 -643 695
rect -701 655 -689 689
rect -655 655 -643 689
rect -701 649 -643 655
rect -509 689 -451 695
rect -509 655 -497 689
rect -463 655 -451 689
rect -509 649 -451 655
rect -317 689 -259 695
rect -317 655 -305 689
rect -271 655 -259 689
rect -317 649 -259 655
rect -125 689 -67 695
rect -125 655 -113 689
rect -79 655 -67 689
rect -125 649 -67 655
rect 67 689 125 695
rect 67 655 79 689
rect 113 655 125 689
rect 67 649 125 655
rect 259 689 317 695
rect 259 655 271 689
rect 305 655 317 689
rect 259 649 317 655
rect 451 689 509 695
rect 451 655 463 689
rect 497 655 509 689
rect 451 649 509 655
rect 643 689 701 695
rect 643 655 655 689
rect 689 655 701 689
rect 643 649 701 655
rect 835 689 893 695
rect 835 655 847 689
rect 881 655 893 689
rect 835 649 893 655
rect 1027 689 1085 695
rect 1027 655 1039 689
rect 1073 655 1085 689
rect 1027 649 1085 655
rect -1085 581 -1027 587
rect -1085 547 -1073 581
rect -1039 547 -1027 581
rect -1085 541 -1027 547
rect -893 581 -835 587
rect -893 547 -881 581
rect -847 547 -835 581
rect -893 541 -835 547
rect -701 581 -643 587
rect -701 547 -689 581
rect -655 547 -643 581
rect -701 541 -643 547
rect -509 581 -451 587
rect -509 547 -497 581
rect -463 547 -451 581
rect -509 541 -451 547
rect -317 581 -259 587
rect -317 547 -305 581
rect -271 547 -259 581
rect -317 541 -259 547
rect -125 581 -67 587
rect -125 547 -113 581
rect -79 547 -67 581
rect -125 541 -67 547
rect 67 581 125 587
rect 67 547 79 581
rect 113 547 125 581
rect 67 541 125 547
rect 259 581 317 587
rect 259 547 271 581
rect 305 547 317 581
rect 259 541 317 547
rect 451 581 509 587
rect 451 547 463 581
rect 497 547 509 581
rect 451 541 509 547
rect 643 581 701 587
rect 643 547 655 581
rect 689 547 701 581
rect 643 541 701 547
rect 835 581 893 587
rect 835 547 847 581
rect 881 547 893 581
rect 835 541 893 547
rect 1027 581 1085 587
rect 1027 547 1039 581
rect 1073 547 1085 581
rect 1027 541 1085 547
rect -1223 497 -1177 509
rect -1223 121 -1217 497
rect -1183 121 -1177 497
rect -1223 109 -1177 121
rect -1127 497 -1081 509
rect -1127 121 -1121 497
rect -1087 121 -1081 497
rect -1127 109 -1081 121
rect -1031 497 -985 509
rect -1031 121 -1025 497
rect -991 121 -985 497
rect -1031 109 -985 121
rect -935 497 -889 509
rect -935 121 -929 497
rect -895 121 -889 497
rect -935 109 -889 121
rect -839 497 -793 509
rect -839 121 -833 497
rect -799 121 -793 497
rect -839 109 -793 121
rect -743 497 -697 509
rect -743 121 -737 497
rect -703 121 -697 497
rect -743 109 -697 121
rect -647 497 -601 509
rect -647 121 -641 497
rect -607 121 -601 497
rect -647 109 -601 121
rect -551 497 -505 509
rect -551 121 -545 497
rect -511 121 -505 497
rect -551 109 -505 121
rect -455 497 -409 509
rect -455 121 -449 497
rect -415 121 -409 497
rect -455 109 -409 121
rect -359 497 -313 509
rect -359 121 -353 497
rect -319 121 -313 497
rect -359 109 -313 121
rect -263 497 -217 509
rect -263 121 -257 497
rect -223 121 -217 497
rect -263 109 -217 121
rect -167 497 -121 509
rect -167 121 -161 497
rect -127 121 -121 497
rect -167 109 -121 121
rect -71 497 -25 509
rect -71 121 -65 497
rect -31 121 -25 497
rect -71 109 -25 121
rect 25 497 71 509
rect 25 121 31 497
rect 65 121 71 497
rect 25 109 71 121
rect 121 497 167 509
rect 121 121 127 497
rect 161 121 167 497
rect 121 109 167 121
rect 217 497 263 509
rect 217 121 223 497
rect 257 121 263 497
rect 217 109 263 121
rect 313 497 359 509
rect 313 121 319 497
rect 353 121 359 497
rect 313 109 359 121
rect 409 497 455 509
rect 409 121 415 497
rect 449 121 455 497
rect 409 109 455 121
rect 505 497 551 509
rect 505 121 511 497
rect 545 121 551 497
rect 505 109 551 121
rect 601 497 647 509
rect 601 121 607 497
rect 641 121 647 497
rect 601 109 647 121
rect 697 497 743 509
rect 697 121 703 497
rect 737 121 743 497
rect 697 109 743 121
rect 793 497 839 509
rect 793 121 799 497
rect 833 121 839 497
rect 793 109 839 121
rect 889 497 935 509
rect 889 121 895 497
rect 929 121 935 497
rect 889 109 935 121
rect 985 497 1031 509
rect 985 121 991 497
rect 1025 121 1031 497
rect 985 109 1031 121
rect 1081 497 1127 509
rect 1081 121 1087 497
rect 1121 121 1127 497
rect 1081 109 1127 121
rect 1177 497 1223 509
rect 1177 121 1183 497
rect 1217 121 1223 497
rect 1177 109 1223 121
rect -1181 71 -1123 77
rect -1181 37 -1169 71
rect -1135 37 -1123 71
rect -1181 31 -1123 37
rect -989 71 -931 77
rect -989 37 -977 71
rect -943 37 -931 71
rect -989 31 -931 37
rect -797 71 -739 77
rect -797 37 -785 71
rect -751 37 -739 71
rect -797 31 -739 37
rect -605 71 -547 77
rect -605 37 -593 71
rect -559 37 -547 71
rect -605 31 -547 37
rect -413 71 -355 77
rect -413 37 -401 71
rect -367 37 -355 71
rect -413 31 -355 37
rect -221 71 -163 77
rect -221 37 -209 71
rect -175 37 -163 71
rect -221 31 -163 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 163 71 221 77
rect 163 37 175 71
rect 209 37 221 71
rect 163 31 221 37
rect 355 71 413 77
rect 355 37 367 71
rect 401 37 413 71
rect 355 31 413 37
rect 547 71 605 77
rect 547 37 559 71
rect 593 37 605 71
rect 547 31 605 37
rect 739 71 797 77
rect 739 37 751 71
rect 785 37 797 71
rect 739 31 797 37
rect 931 71 989 77
rect 931 37 943 71
rect 977 37 989 71
rect 931 31 989 37
rect 1123 71 1181 77
rect 1123 37 1135 71
rect 1169 37 1181 71
rect 1123 31 1181 37
rect -1181 -37 -1123 -31
rect -1181 -71 -1169 -37
rect -1135 -71 -1123 -37
rect -1181 -77 -1123 -71
rect -989 -37 -931 -31
rect -989 -71 -977 -37
rect -943 -71 -931 -37
rect -989 -77 -931 -71
rect -797 -37 -739 -31
rect -797 -71 -785 -37
rect -751 -71 -739 -37
rect -797 -77 -739 -71
rect -605 -37 -547 -31
rect -605 -71 -593 -37
rect -559 -71 -547 -37
rect -605 -77 -547 -71
rect -413 -37 -355 -31
rect -413 -71 -401 -37
rect -367 -71 -355 -37
rect -413 -77 -355 -71
rect -221 -37 -163 -31
rect -221 -71 -209 -37
rect -175 -71 -163 -37
rect -221 -77 -163 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 163 -37 221 -31
rect 163 -71 175 -37
rect 209 -71 221 -37
rect 163 -77 221 -71
rect 355 -37 413 -31
rect 355 -71 367 -37
rect 401 -71 413 -37
rect 355 -77 413 -71
rect 547 -37 605 -31
rect 547 -71 559 -37
rect 593 -71 605 -37
rect 547 -77 605 -71
rect 739 -37 797 -31
rect 739 -71 751 -37
rect 785 -71 797 -37
rect 739 -77 797 -71
rect 931 -37 989 -31
rect 931 -71 943 -37
rect 977 -71 989 -37
rect 931 -77 989 -71
rect 1123 -37 1181 -31
rect 1123 -71 1135 -37
rect 1169 -71 1181 -37
rect 1123 -77 1181 -71
rect -1223 -121 -1177 -109
rect -1223 -497 -1217 -121
rect -1183 -497 -1177 -121
rect -1223 -509 -1177 -497
rect -1127 -121 -1081 -109
rect -1127 -497 -1121 -121
rect -1087 -497 -1081 -121
rect -1127 -509 -1081 -497
rect -1031 -121 -985 -109
rect -1031 -497 -1025 -121
rect -991 -497 -985 -121
rect -1031 -509 -985 -497
rect -935 -121 -889 -109
rect -935 -497 -929 -121
rect -895 -497 -889 -121
rect -935 -509 -889 -497
rect -839 -121 -793 -109
rect -839 -497 -833 -121
rect -799 -497 -793 -121
rect -839 -509 -793 -497
rect -743 -121 -697 -109
rect -743 -497 -737 -121
rect -703 -497 -697 -121
rect -743 -509 -697 -497
rect -647 -121 -601 -109
rect -647 -497 -641 -121
rect -607 -497 -601 -121
rect -647 -509 -601 -497
rect -551 -121 -505 -109
rect -551 -497 -545 -121
rect -511 -497 -505 -121
rect -551 -509 -505 -497
rect -455 -121 -409 -109
rect -455 -497 -449 -121
rect -415 -497 -409 -121
rect -455 -509 -409 -497
rect -359 -121 -313 -109
rect -359 -497 -353 -121
rect -319 -497 -313 -121
rect -359 -509 -313 -497
rect -263 -121 -217 -109
rect -263 -497 -257 -121
rect -223 -497 -217 -121
rect -263 -509 -217 -497
rect -167 -121 -121 -109
rect -167 -497 -161 -121
rect -127 -497 -121 -121
rect -167 -509 -121 -497
rect -71 -121 -25 -109
rect -71 -497 -65 -121
rect -31 -497 -25 -121
rect -71 -509 -25 -497
rect 25 -121 71 -109
rect 25 -497 31 -121
rect 65 -497 71 -121
rect 25 -509 71 -497
rect 121 -121 167 -109
rect 121 -497 127 -121
rect 161 -497 167 -121
rect 121 -509 167 -497
rect 217 -121 263 -109
rect 217 -497 223 -121
rect 257 -497 263 -121
rect 217 -509 263 -497
rect 313 -121 359 -109
rect 313 -497 319 -121
rect 353 -497 359 -121
rect 313 -509 359 -497
rect 409 -121 455 -109
rect 409 -497 415 -121
rect 449 -497 455 -121
rect 409 -509 455 -497
rect 505 -121 551 -109
rect 505 -497 511 -121
rect 545 -497 551 -121
rect 505 -509 551 -497
rect 601 -121 647 -109
rect 601 -497 607 -121
rect 641 -497 647 -121
rect 601 -509 647 -497
rect 697 -121 743 -109
rect 697 -497 703 -121
rect 737 -497 743 -121
rect 697 -509 743 -497
rect 793 -121 839 -109
rect 793 -497 799 -121
rect 833 -497 839 -121
rect 793 -509 839 -497
rect 889 -121 935 -109
rect 889 -497 895 -121
rect 929 -497 935 -121
rect 889 -509 935 -497
rect 985 -121 1031 -109
rect 985 -497 991 -121
rect 1025 -497 1031 -121
rect 985 -509 1031 -497
rect 1081 -121 1127 -109
rect 1081 -497 1087 -121
rect 1121 -497 1127 -121
rect 1081 -509 1127 -497
rect 1177 -121 1223 -109
rect 1177 -497 1183 -121
rect 1217 -497 1223 -121
rect 1177 -509 1223 -497
rect -1085 -547 -1027 -541
rect -1085 -581 -1073 -547
rect -1039 -581 -1027 -547
rect -1085 -587 -1027 -581
rect -893 -547 -835 -541
rect -893 -581 -881 -547
rect -847 -581 -835 -547
rect -893 -587 -835 -581
rect -701 -547 -643 -541
rect -701 -581 -689 -547
rect -655 -581 -643 -547
rect -701 -587 -643 -581
rect -509 -547 -451 -541
rect -509 -581 -497 -547
rect -463 -581 -451 -547
rect -509 -587 -451 -581
rect -317 -547 -259 -541
rect -317 -581 -305 -547
rect -271 -581 -259 -547
rect -317 -587 -259 -581
rect -125 -547 -67 -541
rect -125 -581 -113 -547
rect -79 -581 -67 -547
rect -125 -587 -67 -581
rect 67 -547 125 -541
rect 67 -581 79 -547
rect 113 -581 125 -547
rect 67 -587 125 -581
rect 259 -547 317 -541
rect 259 -581 271 -547
rect 305 -581 317 -547
rect 259 -587 317 -581
rect 451 -547 509 -541
rect 451 -581 463 -547
rect 497 -581 509 -547
rect 451 -587 509 -581
rect 643 -547 701 -541
rect 643 -581 655 -547
rect 689 -581 701 -547
rect 643 -587 701 -581
rect 835 -547 893 -541
rect 835 -581 847 -547
rect 881 -581 893 -547
rect 835 -587 893 -581
rect 1027 -547 1085 -541
rect 1027 -581 1039 -547
rect 1073 -581 1085 -547
rect 1027 -587 1085 -581
rect -1085 -655 -1027 -649
rect -1085 -689 -1073 -655
rect -1039 -689 -1027 -655
rect -1085 -695 -1027 -689
rect -893 -655 -835 -649
rect -893 -689 -881 -655
rect -847 -689 -835 -655
rect -893 -695 -835 -689
rect -701 -655 -643 -649
rect -701 -689 -689 -655
rect -655 -689 -643 -655
rect -701 -695 -643 -689
rect -509 -655 -451 -649
rect -509 -689 -497 -655
rect -463 -689 -451 -655
rect -509 -695 -451 -689
rect -317 -655 -259 -649
rect -317 -689 -305 -655
rect -271 -689 -259 -655
rect -317 -695 -259 -689
rect -125 -655 -67 -649
rect -125 -689 -113 -655
rect -79 -689 -67 -655
rect -125 -695 -67 -689
rect 67 -655 125 -649
rect 67 -689 79 -655
rect 113 -689 125 -655
rect 67 -695 125 -689
rect 259 -655 317 -649
rect 259 -689 271 -655
rect 305 -689 317 -655
rect 259 -695 317 -689
rect 451 -655 509 -649
rect 451 -689 463 -655
rect 497 -689 509 -655
rect 451 -695 509 -689
rect 643 -655 701 -649
rect 643 -689 655 -655
rect 689 -689 701 -655
rect 643 -695 701 -689
rect 835 -655 893 -649
rect 835 -689 847 -655
rect 881 -689 893 -655
rect 835 -695 893 -689
rect 1027 -655 1085 -649
rect 1027 -689 1039 -655
rect 1073 -689 1085 -655
rect 1027 -695 1085 -689
rect -1223 -739 -1177 -727
rect -1223 -1115 -1217 -739
rect -1183 -1115 -1177 -739
rect -1223 -1127 -1177 -1115
rect -1127 -739 -1081 -727
rect -1127 -1115 -1121 -739
rect -1087 -1115 -1081 -739
rect -1127 -1127 -1081 -1115
rect -1031 -739 -985 -727
rect -1031 -1115 -1025 -739
rect -991 -1115 -985 -739
rect -1031 -1127 -985 -1115
rect -935 -739 -889 -727
rect -935 -1115 -929 -739
rect -895 -1115 -889 -739
rect -935 -1127 -889 -1115
rect -839 -739 -793 -727
rect -839 -1115 -833 -739
rect -799 -1115 -793 -739
rect -839 -1127 -793 -1115
rect -743 -739 -697 -727
rect -743 -1115 -737 -739
rect -703 -1115 -697 -739
rect -743 -1127 -697 -1115
rect -647 -739 -601 -727
rect -647 -1115 -641 -739
rect -607 -1115 -601 -739
rect -647 -1127 -601 -1115
rect -551 -739 -505 -727
rect -551 -1115 -545 -739
rect -511 -1115 -505 -739
rect -551 -1127 -505 -1115
rect -455 -739 -409 -727
rect -455 -1115 -449 -739
rect -415 -1115 -409 -739
rect -455 -1127 -409 -1115
rect -359 -739 -313 -727
rect -359 -1115 -353 -739
rect -319 -1115 -313 -739
rect -359 -1127 -313 -1115
rect -263 -739 -217 -727
rect -263 -1115 -257 -739
rect -223 -1115 -217 -739
rect -263 -1127 -217 -1115
rect -167 -739 -121 -727
rect -167 -1115 -161 -739
rect -127 -1115 -121 -739
rect -167 -1127 -121 -1115
rect -71 -739 -25 -727
rect -71 -1115 -65 -739
rect -31 -1115 -25 -739
rect -71 -1127 -25 -1115
rect 25 -739 71 -727
rect 25 -1115 31 -739
rect 65 -1115 71 -739
rect 25 -1127 71 -1115
rect 121 -739 167 -727
rect 121 -1115 127 -739
rect 161 -1115 167 -739
rect 121 -1127 167 -1115
rect 217 -739 263 -727
rect 217 -1115 223 -739
rect 257 -1115 263 -739
rect 217 -1127 263 -1115
rect 313 -739 359 -727
rect 313 -1115 319 -739
rect 353 -1115 359 -739
rect 313 -1127 359 -1115
rect 409 -739 455 -727
rect 409 -1115 415 -739
rect 449 -1115 455 -739
rect 409 -1127 455 -1115
rect 505 -739 551 -727
rect 505 -1115 511 -739
rect 545 -1115 551 -739
rect 505 -1127 551 -1115
rect 601 -739 647 -727
rect 601 -1115 607 -739
rect 641 -1115 647 -739
rect 601 -1127 647 -1115
rect 697 -739 743 -727
rect 697 -1115 703 -739
rect 737 -1115 743 -739
rect 697 -1127 743 -1115
rect 793 -739 839 -727
rect 793 -1115 799 -739
rect 833 -1115 839 -739
rect 793 -1127 839 -1115
rect 889 -739 935 -727
rect 889 -1115 895 -739
rect 929 -1115 935 -739
rect 889 -1127 935 -1115
rect 985 -739 1031 -727
rect 985 -1115 991 -739
rect 1025 -1115 1031 -739
rect 985 -1127 1031 -1115
rect 1081 -739 1127 -727
rect 1081 -1115 1087 -739
rect 1121 -1115 1127 -739
rect 1081 -1127 1127 -1115
rect 1177 -739 1223 -727
rect 1177 -1115 1183 -739
rect 1217 -1115 1223 -739
rect 1177 -1127 1223 -1115
rect -1181 -1165 -1123 -1159
rect -1181 -1199 -1169 -1165
rect -1135 -1199 -1123 -1165
rect -1181 -1205 -1123 -1199
rect -989 -1165 -931 -1159
rect -989 -1199 -977 -1165
rect -943 -1199 -931 -1165
rect -989 -1205 -931 -1199
rect -797 -1165 -739 -1159
rect -797 -1199 -785 -1165
rect -751 -1199 -739 -1165
rect -797 -1205 -739 -1199
rect -605 -1165 -547 -1159
rect -605 -1199 -593 -1165
rect -559 -1199 -547 -1165
rect -605 -1205 -547 -1199
rect -413 -1165 -355 -1159
rect -413 -1199 -401 -1165
rect -367 -1199 -355 -1165
rect -413 -1205 -355 -1199
rect -221 -1165 -163 -1159
rect -221 -1199 -209 -1165
rect -175 -1199 -163 -1165
rect -221 -1205 -163 -1199
rect -29 -1165 29 -1159
rect -29 -1199 -17 -1165
rect 17 -1199 29 -1165
rect -29 -1205 29 -1199
rect 163 -1165 221 -1159
rect 163 -1199 175 -1165
rect 209 -1199 221 -1165
rect 163 -1205 221 -1199
rect 355 -1165 413 -1159
rect 355 -1199 367 -1165
rect 401 -1199 413 -1165
rect 355 -1205 413 -1199
rect 547 -1165 605 -1159
rect 547 -1199 559 -1165
rect 593 -1199 605 -1165
rect 547 -1205 605 -1199
rect 739 -1165 797 -1159
rect 739 -1199 751 -1165
rect 785 -1199 797 -1165
rect 739 -1205 797 -1199
rect 931 -1165 989 -1159
rect 931 -1199 943 -1165
rect 977 -1199 989 -1165
rect 931 -1205 989 -1199
rect 1123 -1165 1181 -1159
rect 1123 -1199 1135 -1165
rect 1169 -1199 1181 -1165
rect 1123 -1205 1181 -1199
<< properties >>
string FIXED_BBOX -1314 -1284 1314 1284
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 4 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
