magic
tech sky130A
magscale 1 2
timestamp 1646060485
<< metal3 >>
rect -1350 1572 1349 1600
rect -1350 -1572 1265 1572
rect 1329 -1572 1349 1572
rect -1350 -1600 1349 -1572
<< via3 >>
rect 1265 -1572 1329 1572
<< mimcap >>
rect -1250 1460 1150 1500
rect -1250 -1460 -1210 1460
rect 1110 -1460 1150 1460
rect -1250 -1500 1150 -1460
<< mimcapcontact >>
rect -1210 -1460 1110 1460
<< metal4 >>
rect 1249 1572 1345 1588
rect -1211 1460 1111 1461
rect -1211 -1460 -1210 1460
rect 1110 -1460 1111 1460
rect -1211 -1461 1111 -1460
rect 1249 -1572 1265 1572
rect 1329 -1572 1345 1572
rect 1249 -1588 1345 -1572
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -1350 -1600 1250 1600
string parameters w 12 l 15 val 370.26 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
