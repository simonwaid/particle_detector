magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< nwell >>
rect 122 3370 1488 3436
rect 122 2852 1488 2898
rect 112 640 1234 706
rect 130 634 160 640
rect 322 634 352 640
rect 514 634 544 640
rect 706 634 736 640
rect 898 634 928 640
rect 1090 634 1120 640
rect 226 178 256 184
rect 418 178 448 184
rect 610 178 640 184
rect 802 178 832 184
rect 994 178 1024 184
rect 1186 178 1216 184
rect 112 112 1234 178
<< poly >>
rect 122 4006 1488 4072
rect 122 3488 1488 3534
rect 122 3370 1488 3436
rect 122 2852 1488 2898
rect 112 2598 1234 2614
rect 112 2564 224 2598
rect 258 2564 416 2598
rect 450 2564 608 2598
rect 642 2564 800 2598
rect 834 2564 992 2598
rect 1026 2564 1184 2598
rect 1218 2564 1234 2598
rect 112 2548 1234 2564
rect 226 2542 256 2548
rect 418 2542 448 2548
rect 610 2542 640 2548
rect 802 2542 832 2548
rect 994 2542 1024 2548
rect 1186 2542 1216 2548
rect 130 2086 160 2092
rect 322 2086 352 2092
rect 514 2086 544 2092
rect 706 2086 736 2092
rect 898 2086 928 2092
rect 1090 2086 1120 2092
rect 112 2070 1234 2086
rect 112 2036 128 2070
rect 162 2036 320 2070
rect 354 2036 512 2070
rect 546 2036 704 2070
rect 738 2036 896 2070
rect 930 2036 1088 2070
rect 1122 2036 1234 2070
rect 112 2020 1234 2036
rect 112 1962 1234 1978
rect 112 1928 128 1962
rect 162 1928 320 1962
rect 354 1928 512 1962
rect 546 1928 704 1962
rect 738 1928 896 1962
rect 930 1928 1088 1962
rect 1122 1928 1234 1962
rect 112 1912 1234 1928
rect 130 1906 160 1912
rect 322 1906 352 1912
rect 514 1906 544 1912
rect 706 1906 736 1912
rect 898 1906 928 1912
rect 1090 1906 1120 1912
rect 226 1450 256 1456
rect 418 1450 448 1456
rect 610 1450 640 1456
rect 802 1450 832 1456
rect 994 1450 1024 1456
rect 1186 1450 1216 1456
rect 112 1434 1234 1450
rect 112 1400 224 1434
rect 258 1400 416 1434
rect 450 1400 608 1434
rect 642 1400 800 1434
rect 834 1400 992 1434
rect 1026 1400 1184 1434
rect 1218 1400 1234 1434
rect 112 1384 1234 1400
rect 112 1326 1234 1342
rect 112 1292 224 1326
rect 258 1292 416 1326
rect 450 1292 608 1326
rect 642 1292 800 1326
rect 834 1292 992 1326
rect 1026 1292 1184 1326
rect 1218 1292 1234 1326
rect 112 1276 1234 1292
rect 226 1270 256 1276
rect 418 1270 448 1276
rect 610 1270 640 1276
rect 802 1270 832 1276
rect 994 1270 1024 1276
rect 1186 1270 1216 1276
rect 130 814 160 820
rect 322 814 352 820
rect 514 814 544 820
rect 706 814 736 820
rect 898 814 928 820
rect 1090 814 1120 820
rect 112 798 1234 814
rect 112 764 128 798
rect 162 764 320 798
rect 354 764 512 798
rect 546 764 704 798
rect 738 764 896 798
rect 930 764 1088 798
rect 1122 764 1234 798
rect 112 748 1234 764
rect 112 690 1234 706
rect 112 656 128 690
rect 162 656 320 690
rect 354 656 512 690
rect 546 656 704 690
rect 738 656 896 690
rect 930 656 1088 690
rect 1122 656 1234 690
rect 112 640 1234 656
rect 130 634 160 640
rect 322 634 352 640
rect 514 634 544 640
rect 706 634 736 640
rect 898 634 928 640
rect 1090 634 1120 640
rect 226 178 256 184
rect 418 178 448 184
rect 610 178 640 184
rect 802 178 832 184
rect 994 178 1024 184
rect 1186 178 1216 184
rect 112 162 1234 178
rect 112 128 224 162
rect 258 128 416 162
rect 450 128 608 162
rect 642 128 800 162
rect 834 128 992 162
rect 1026 128 1184 162
rect 1218 128 1234 162
rect 112 112 1234 128
<< polycont >>
rect 224 2564 258 2598
rect 416 2564 450 2598
rect 608 2564 642 2598
rect 800 2564 834 2598
rect 992 2564 1026 2598
rect 1184 2564 1218 2598
rect 128 2036 162 2070
rect 320 2036 354 2070
rect 512 2036 546 2070
rect 704 2036 738 2070
rect 896 2036 930 2070
rect 1088 2036 1122 2070
rect 128 1928 162 1962
rect 320 1928 354 1962
rect 512 1928 546 1962
rect 704 1928 738 1962
rect 896 1928 930 1962
rect 1088 1928 1122 1962
rect 224 1400 258 1434
rect 416 1400 450 1434
rect 608 1400 642 1434
rect 800 1400 834 1434
rect 992 1400 1026 1434
rect 1184 1400 1218 1434
rect 224 1292 258 1326
rect 416 1292 450 1326
rect 608 1292 642 1326
rect 800 1292 834 1326
rect 992 1292 1026 1326
rect 1184 1292 1218 1326
rect 128 764 162 798
rect 320 764 354 798
rect 512 764 546 798
rect 704 764 738 798
rect 896 764 930 798
rect 1088 764 1122 798
rect 128 656 162 690
rect 320 656 354 690
rect 512 656 546 690
rect 704 656 738 690
rect 896 656 930 690
rect 1088 656 1122 690
rect 224 128 258 162
rect 416 128 450 162
rect 608 128 642 162
rect 800 128 834 162
rect 992 128 1026 162
rect 1184 128 1218 162
<< locali >>
rect 122 4022 1488 4056
rect 122 3494 1488 3528
rect 122 3386 1488 3420
rect 1590 3350 1630 4140
rect 122 2858 1488 2892
rect 1590 2780 1630 3210
rect 1360 2770 1630 2780
rect -30 2760 1630 2770
rect -30 2690 1590 2760
rect 112 2564 224 2598
rect 258 2564 416 2598
rect 450 2564 608 2598
rect 642 2564 800 2598
rect 834 2564 992 2598
rect 1026 2564 1184 2598
rect 1218 2564 1234 2598
rect 112 2036 128 2070
rect 162 2036 320 2070
rect 354 2036 512 2070
rect 546 2036 704 2070
rect 738 2036 896 2070
rect 930 2036 1088 2070
rect 1122 2036 1234 2070
rect 112 1928 128 1962
rect 162 1928 320 1962
rect 354 1928 512 1962
rect 546 1928 704 1962
rect 738 1928 896 1962
rect 930 1928 1088 1962
rect 1122 1928 1234 1962
rect 112 1400 224 1434
rect 258 1400 416 1434
rect 450 1400 608 1434
rect 642 1400 800 1434
rect 834 1400 992 1434
rect 1026 1400 1184 1434
rect 1218 1400 1234 1434
rect 112 1292 224 1326
rect 258 1292 416 1326
rect 450 1292 608 1326
rect 642 1292 800 1326
rect 834 1292 992 1326
rect 1026 1292 1184 1326
rect 1218 1292 1234 1326
rect 112 764 128 798
rect 162 764 320 798
rect 354 764 512 798
rect 546 764 704 798
rect 738 764 896 798
rect 930 764 1088 798
rect 1122 764 1234 798
rect 112 656 128 690
rect 162 656 320 690
rect 354 656 512 690
rect 546 656 704 690
rect 738 656 896 690
rect 930 656 1088 690
rect 1122 656 1234 690
rect 112 128 224 162
rect 258 128 416 162
rect 450 128 608 162
rect 642 128 800 162
rect 834 128 992 162
rect 1026 128 1184 162
rect 1218 128 1234 162
rect 1360 30 1590 2690
<< viali >>
rect 1590 3210 1650 3350
rect 224 2564 258 2598
rect 416 2564 450 2598
rect 608 2564 642 2598
rect 800 2564 834 2598
rect 992 2564 1026 2598
rect 1184 2564 1218 2598
rect 128 2036 162 2070
rect 320 2036 354 2070
rect 512 2036 546 2070
rect 704 2036 738 2070
rect 896 2036 930 2070
rect 1088 2036 1122 2070
rect 128 1928 162 1962
rect 320 1928 354 1962
rect 512 1928 546 1962
rect 704 1928 738 1962
rect 896 1928 930 1962
rect 1088 1928 1122 1962
rect 224 1400 258 1434
rect 416 1400 450 1434
rect 608 1400 642 1434
rect 800 1400 834 1434
rect 992 1400 1026 1434
rect 1184 1400 1218 1434
rect 224 1292 258 1326
rect 416 1292 450 1326
rect 608 1292 642 1326
rect 800 1292 834 1326
rect 992 1292 1026 1326
rect 1184 1292 1218 1326
rect 128 764 162 798
rect 320 764 354 798
rect 512 764 546 798
rect 704 764 738 798
rect 896 764 930 798
rect 1088 764 1122 798
rect 128 656 162 690
rect 320 656 354 690
rect 512 656 546 690
rect 704 656 738 690
rect 896 656 930 690
rect 1088 656 1122 690
rect 224 128 258 162
rect 416 128 450 162
rect 608 128 642 162
rect 800 128 834 162
rect 992 128 1026 162
rect 1184 128 1218 162
<< metal1 >>
rect -30 4010 1490 4070
rect -30 3540 20 4010
rect 178 3800 188 3976
rect 242 3800 252 3976
rect 414 3800 424 3976
rect 478 3800 488 3976
rect 650 3800 660 3976
rect 714 3800 724 3976
rect 886 3800 896 3976
rect 950 3800 960 3976
rect 1122 3800 1132 3976
rect 1186 3800 1196 3976
rect 1358 3800 1368 3976
rect 1422 3800 1432 3976
rect 60 3574 70 3750
rect 124 3574 134 3750
rect 296 3574 306 3750
rect 360 3574 370 3750
rect 532 3574 542 3750
rect 596 3574 606 3750
rect 768 3574 778 3750
rect 832 3574 842 3750
rect 1004 3574 1014 3750
rect 1068 3574 1078 3750
rect 1240 3574 1250 3750
rect 1304 3574 1314 3750
rect 1476 3574 1486 3750
rect 1540 3574 1550 3750
rect -30 3480 1490 3540
rect -30 3440 20 3480
rect -30 3380 1490 3440
rect -30 2900 20 3380
rect 1584 3350 1656 3362
rect 178 3164 188 3340
rect 242 3164 252 3340
rect 414 3164 424 3340
rect 478 3164 488 3340
rect 650 3164 660 3340
rect 714 3164 724 3340
rect 886 3164 896 3340
rect 950 3164 960 3340
rect 1122 3164 1132 3340
rect 1186 3164 1196 3340
rect 1358 3164 1368 3340
rect 1422 3164 1432 3340
rect 1580 3210 1590 3350
rect 1650 3210 1660 3350
rect 1584 3198 1656 3210
rect 60 2938 70 3114
rect 124 2938 134 3114
rect 296 2938 306 3114
rect 360 2938 370 3114
rect 532 2938 542 3114
rect 596 2938 606 3114
rect 768 2938 778 3114
rect 832 2938 842 3114
rect 1004 2938 1014 3114
rect 1068 2938 1078 3114
rect 1240 2938 1250 3114
rect 1304 2938 1314 3114
rect 1476 2938 1486 3114
rect 1540 2938 1550 3114
rect -30 2840 1490 2900
rect -30 2610 20 2840
rect -30 2598 1310 2610
rect -30 2564 224 2598
rect 258 2564 416 2598
rect 450 2564 608 2598
rect 642 2564 800 2598
rect 834 2564 992 2598
rect 1026 2564 1184 2598
rect 1218 2564 1310 2598
rect -30 2550 1310 2564
rect -30 2080 20 2550
rect 60 2342 70 2518
rect 124 2342 134 2518
rect 252 2342 262 2518
rect 316 2342 326 2518
rect 444 2342 454 2518
rect 508 2342 518 2518
rect 636 2342 646 2518
rect 700 2342 710 2518
rect 828 2342 838 2518
rect 892 2342 902 2518
rect 1020 2342 1030 2518
rect 1084 2342 1094 2518
rect 1212 2342 1222 2518
rect 1276 2342 1286 2518
rect 156 2116 166 2292
rect 220 2116 230 2292
rect 348 2116 358 2292
rect 412 2116 422 2292
rect 540 2116 550 2292
rect 604 2116 614 2292
rect 732 2116 742 2292
rect 796 2116 806 2292
rect 924 2116 934 2292
rect 988 2116 998 2292
rect 1116 2116 1126 2292
rect 1180 2116 1190 2292
rect -30 2070 1310 2080
rect -30 2036 128 2070
rect 162 2036 320 2070
rect 354 2036 512 2070
rect 546 2036 704 2070
rect 738 2036 896 2070
rect 930 2036 1088 2070
rect 1122 2036 1310 2070
rect -30 2020 1310 2036
rect -30 1980 20 2020
rect -30 1962 1310 1980
rect -30 1928 128 1962
rect 162 1928 320 1962
rect 354 1928 512 1962
rect 546 1928 704 1962
rect 738 1928 896 1962
rect 930 1928 1088 1962
rect 1122 1928 1310 1962
rect -30 1920 1310 1928
rect -30 1440 20 1920
rect 156 1706 166 1882
rect 220 1706 230 1882
rect 348 1706 358 1882
rect 412 1706 422 1882
rect 540 1706 550 1882
rect 604 1706 614 1882
rect 732 1706 742 1882
rect 796 1706 806 1882
rect 924 1706 934 1882
rect 988 1706 998 1882
rect 1116 1706 1126 1882
rect 1180 1706 1190 1882
rect 60 1480 70 1656
rect 124 1480 134 1656
rect 252 1480 262 1656
rect 316 1480 326 1656
rect 444 1480 454 1656
rect 508 1480 518 1656
rect 636 1480 646 1656
rect 700 1480 710 1656
rect 828 1480 838 1656
rect 892 1480 902 1656
rect 1020 1480 1030 1656
rect 1084 1480 1094 1656
rect 1212 1480 1222 1656
rect 1276 1480 1286 1656
rect -30 1434 1310 1440
rect -30 1400 224 1434
rect 258 1400 416 1434
rect 450 1400 608 1434
rect 642 1400 800 1434
rect 834 1400 992 1434
rect 1026 1400 1184 1434
rect 1218 1400 1310 1434
rect -30 1380 1310 1400
rect -30 1340 20 1380
rect -30 1326 1310 1340
rect -30 1292 224 1326
rect 258 1292 416 1326
rect 450 1292 608 1326
rect 642 1292 800 1326
rect 834 1292 992 1326
rect 1026 1292 1184 1326
rect 1218 1292 1310 1326
rect -30 1280 1310 1292
rect -30 810 20 1280
rect 60 1070 70 1246
rect 124 1070 134 1246
rect 252 1070 262 1246
rect 316 1070 326 1246
rect 444 1070 454 1246
rect 508 1070 518 1246
rect 636 1070 646 1246
rect 700 1070 710 1246
rect 828 1070 838 1246
rect 892 1070 902 1246
rect 1020 1070 1030 1246
rect 1084 1070 1094 1246
rect 1212 1070 1222 1246
rect 1276 1070 1286 1246
rect 156 844 166 1020
rect 220 844 230 1020
rect 348 844 358 1020
rect 412 844 422 1020
rect 540 844 550 1020
rect 604 844 614 1020
rect 732 844 742 1020
rect 796 844 806 1020
rect 924 844 934 1020
rect 988 844 998 1020
rect 1116 844 1126 1020
rect 1180 844 1190 1020
rect -30 798 1310 810
rect -30 764 128 798
rect 162 764 320 798
rect 354 764 512 798
rect 546 764 704 798
rect 738 764 896 798
rect 930 764 1088 798
rect 1122 764 1310 798
rect -30 750 1310 764
rect -30 710 20 750
rect -30 690 1310 710
rect -30 656 128 690
rect 162 656 320 690
rect 354 656 512 690
rect 546 656 704 690
rect 738 656 896 690
rect 930 656 1088 690
rect 1122 656 1310 690
rect -30 650 1310 656
rect -30 170 20 650
rect 156 434 166 610
rect 220 434 230 610
rect 348 434 358 610
rect 412 434 422 610
rect 540 434 550 610
rect 604 434 614 610
rect 732 434 742 610
rect 796 434 806 610
rect 924 434 934 610
rect 988 434 998 610
rect 1116 434 1126 610
rect 1180 434 1190 610
rect 60 208 70 384
rect 124 208 134 384
rect 252 208 262 384
rect 316 208 326 384
rect 444 208 454 384
rect 508 208 518 384
rect 636 208 646 384
rect 700 208 710 384
rect 828 208 838 384
rect 892 208 902 384
rect 1020 208 1030 384
rect 1084 208 1094 384
rect 1212 208 1222 384
rect 1276 208 1286 384
rect -30 162 1310 170
rect -30 128 224 162
rect 258 128 416 162
rect 450 128 608 162
rect 642 128 800 162
rect 834 128 992 162
rect 1026 128 1184 162
rect 1218 128 1310 162
rect -30 110 1310 128
<< via1 >>
rect 188 3800 242 3976
rect 424 3800 478 3976
rect 660 3800 714 3976
rect 896 3800 950 3976
rect 1132 3800 1186 3976
rect 1368 3800 1422 3976
rect 70 3574 124 3750
rect 306 3574 360 3750
rect 542 3574 596 3750
rect 778 3574 832 3750
rect 1014 3574 1068 3750
rect 1250 3574 1304 3750
rect 1486 3574 1540 3750
rect 188 3164 242 3340
rect 424 3164 478 3340
rect 660 3164 714 3340
rect 896 3164 950 3340
rect 1132 3164 1186 3340
rect 1368 3164 1422 3340
rect 1590 3210 1650 3350
rect 70 2938 124 3114
rect 306 2938 360 3114
rect 542 2938 596 3114
rect 778 2938 832 3114
rect 1014 2938 1068 3114
rect 1250 2938 1304 3114
rect 1486 2938 1540 3114
rect 70 2342 124 2518
rect 262 2342 316 2518
rect 454 2342 508 2518
rect 646 2342 700 2518
rect 838 2342 892 2518
rect 1030 2342 1084 2518
rect 1222 2342 1276 2518
rect 166 2116 220 2292
rect 358 2116 412 2292
rect 550 2116 604 2292
rect 742 2116 796 2292
rect 934 2116 988 2292
rect 1126 2116 1180 2292
rect 166 1706 220 1882
rect 358 1706 412 1882
rect 550 1706 604 1882
rect 742 1706 796 1882
rect 934 1706 988 1882
rect 1126 1706 1180 1882
rect 70 1480 124 1656
rect 262 1480 316 1656
rect 454 1480 508 1656
rect 646 1480 700 1656
rect 838 1480 892 1656
rect 1030 1480 1084 1656
rect 1222 1480 1276 1656
rect 70 1070 124 1246
rect 262 1070 316 1246
rect 454 1070 508 1246
rect 646 1070 700 1246
rect 838 1070 892 1246
rect 1030 1070 1084 1246
rect 1222 1070 1276 1246
rect 166 844 220 1020
rect 358 844 412 1020
rect 550 844 604 1020
rect 742 844 796 1020
rect 934 844 988 1020
rect 1126 844 1180 1020
rect 166 434 220 610
rect 358 434 412 610
rect 550 434 604 610
rect 742 434 796 610
rect 934 434 988 610
rect 1126 434 1180 610
rect 70 208 124 384
rect 262 208 316 384
rect 454 208 508 384
rect 646 208 700 384
rect 838 208 892 384
rect 1030 208 1084 384
rect 1222 208 1276 384
<< metal2 >>
rect 0 4160 420 4170
rect 1150 4160 1570 4170
rect 420 3976 1150 3990
rect 420 3840 424 3976
rect 0 3830 188 3840
rect 242 3830 424 3840
rect 188 3790 242 3800
rect 478 3830 660 3976
rect 424 3790 478 3800
rect 714 3830 896 3976
rect 660 3790 714 3800
rect 950 3830 1132 3976
rect 896 3790 950 3800
rect 1186 3830 1368 3840
rect 1132 3790 1186 3800
rect 1422 3830 1570 3840
rect 1368 3790 1422 3800
rect 70 3750 124 3760
rect 60 3574 70 3720
rect 306 3750 360 3760
rect 124 3574 306 3720
rect 542 3750 596 3760
rect 360 3710 542 3720
rect 778 3750 832 3760
rect 596 3710 778 3720
rect 1014 3750 1068 3760
rect 832 3710 1014 3720
rect 1250 3750 1304 3760
rect 360 3574 520 3710
rect 1068 3574 1250 3720
rect 1486 3750 1540 3760
rect 1304 3574 1486 3720
rect 1540 3574 1550 3720
rect 60 3560 520 3574
rect 1040 3560 1550 3574
rect 520 3540 1040 3550
rect 0 3470 420 3480
rect 1150 3470 1570 3480
rect 420 3340 1150 3360
rect 1570 3350 1650 3360
rect 420 3210 424 3340
rect 0 3200 188 3210
rect 242 3200 424 3210
rect 188 3154 242 3164
rect 478 3200 660 3340
rect 424 3154 478 3164
rect 714 3200 896 3340
rect 660 3154 714 3164
rect 950 3200 1132 3340
rect 1570 3210 1590 3350
rect 896 3154 950 3164
rect 1186 3200 1368 3210
rect 1132 3154 1186 3164
rect 1422 3200 1650 3210
rect 1368 3154 1422 3164
rect 70 3114 124 3124
rect 60 2938 70 3080
rect 306 3114 360 3124
rect 124 2938 306 3080
rect 542 3114 596 3124
rect 360 3070 542 3080
rect 778 3114 832 3124
rect 596 3070 778 3080
rect 1014 3114 1068 3124
rect 832 3070 1014 3080
rect 1250 3114 1304 3124
rect 360 2938 520 3070
rect 1068 2938 1250 3080
rect 1486 3114 1540 3124
rect 1304 2938 1486 3080
rect 1540 2938 1550 3080
rect 60 2920 520 2938
rect 1040 2920 1550 2938
rect 520 2900 1040 2910
rect 520 2540 1040 2550
rect 60 2518 520 2530
rect 1040 2518 1280 2530
rect 60 2370 70 2518
rect 124 2370 262 2518
rect 70 2332 124 2342
rect 316 2370 454 2518
rect 262 2332 316 2342
rect 508 2380 520 2518
rect 508 2370 646 2380
rect 454 2332 508 2342
rect 700 2370 838 2380
rect 646 2332 700 2342
rect 892 2370 1030 2380
rect 838 2332 892 2342
rect 1084 2370 1222 2518
rect 1030 2332 1084 2342
rect 1276 2370 1280 2518
rect 1222 2332 1276 2342
rect 166 2292 220 2302
rect 0 2250 166 2260
rect 358 2292 412 2302
rect 220 2250 358 2260
rect 550 2292 604 2302
rect 412 2250 550 2260
rect 420 2116 550 2250
rect 742 2292 796 2302
rect 604 2116 742 2260
rect 934 2292 988 2302
rect 796 2116 934 2260
rect 1126 2292 1180 2302
rect 988 2116 1126 2260
rect 1180 2250 1570 2260
rect 420 1882 1150 2116
rect 420 1750 550 1882
rect 0 1740 166 1750
rect 220 1740 358 1750
rect 166 1696 220 1706
rect 412 1740 550 1750
rect 358 1696 412 1706
rect 604 1740 742 1882
rect 550 1696 604 1706
rect 796 1740 934 1882
rect 742 1696 796 1706
rect 988 1740 1126 1882
rect 934 1696 988 1706
rect 1180 1740 1570 1750
rect 1126 1696 1180 1706
rect 70 1656 124 1666
rect 60 1480 70 1620
rect 262 1656 316 1666
rect 124 1480 262 1620
rect 454 1656 508 1666
rect 316 1480 454 1620
rect 646 1656 700 1666
rect 508 1610 646 1620
rect 838 1656 892 1666
rect 700 1610 838 1620
rect 1030 1656 1084 1666
rect 892 1610 1030 1620
rect 1222 1656 1276 1666
rect 508 1480 520 1610
rect 1084 1480 1222 1620
rect 1276 1480 1280 1620
rect 60 1460 520 1480
rect 1040 1460 1280 1480
rect 520 1440 1040 1450
rect 520 1270 1040 1280
rect 60 1246 520 1260
rect 1040 1246 1280 1260
rect 60 1100 70 1246
rect 124 1100 262 1246
rect 70 1060 124 1070
rect 316 1100 454 1246
rect 262 1060 316 1070
rect 508 1110 520 1246
rect 508 1100 646 1110
rect 454 1060 508 1070
rect 700 1100 838 1110
rect 646 1060 700 1070
rect 892 1100 1030 1110
rect 838 1060 892 1070
rect 1084 1100 1222 1246
rect 1030 1060 1084 1070
rect 1276 1100 1280 1246
rect 1222 1060 1276 1070
rect 166 1020 220 1030
rect 0 980 166 990
rect 358 1020 412 1030
rect 220 980 358 990
rect 550 1020 604 1030
rect 412 980 550 990
rect 420 844 550 980
rect 742 1020 796 1030
rect 604 844 742 990
rect 934 1020 988 1030
rect 796 844 934 990
rect 1126 1020 1180 1030
rect 988 844 1126 990
rect 1180 980 1570 990
rect 420 740 1150 844
rect 0 730 1570 740
rect 520 640 1040 650
rect 160 610 520 630
rect 1040 610 1190 630
rect 160 470 166 610
rect 220 470 358 610
rect 166 424 220 434
rect 412 480 520 610
rect 1040 480 1126 610
rect 412 470 550 480
rect 358 424 412 434
rect 604 470 742 480
rect 550 424 604 434
rect 796 470 934 480
rect 742 424 796 434
rect 988 470 1126 480
rect 934 424 988 434
rect 1180 470 1190 610
rect 1126 424 1180 434
rect 70 384 124 394
rect 0 340 70 350
rect 262 384 316 394
rect 124 340 262 350
rect 454 384 508 394
rect 316 340 454 350
rect 420 208 454 340
rect 646 384 700 394
rect 508 208 646 350
rect 838 384 892 394
rect 700 208 838 350
rect 1030 384 1084 394
rect 892 208 1030 350
rect 1222 384 1276 394
rect 1084 340 1222 350
rect 1276 340 1570 350
rect 1084 208 1150 340
rect 420 100 1150 208
rect 0 90 1570 100
<< via2 >>
rect 0 3976 420 4160
rect 1150 3976 1570 4160
rect 0 3840 188 3976
rect 188 3840 242 3976
rect 242 3840 420 3976
rect 1150 3840 1186 3976
rect 1186 3840 1368 3976
rect 1368 3840 1422 3976
rect 1422 3840 1570 3976
rect 520 3574 542 3710
rect 542 3574 596 3710
rect 596 3574 778 3710
rect 778 3574 832 3710
rect 832 3574 1014 3710
rect 1014 3574 1040 3710
rect 520 3550 1040 3574
rect 0 3340 420 3470
rect 1150 3340 1570 3470
rect 0 3210 188 3340
rect 188 3210 242 3340
rect 242 3210 420 3340
rect 1150 3210 1186 3340
rect 1186 3210 1368 3340
rect 1368 3210 1422 3340
rect 1422 3210 1570 3340
rect 520 2938 542 3070
rect 542 2938 596 3070
rect 596 2938 778 3070
rect 778 2938 832 3070
rect 832 2938 1014 3070
rect 1014 2938 1040 3070
rect 520 2910 1040 2938
rect 520 2518 1040 2540
rect 520 2380 646 2518
rect 646 2380 700 2518
rect 700 2380 838 2518
rect 838 2380 892 2518
rect 892 2380 1030 2518
rect 1030 2380 1040 2518
rect 0 2116 166 2250
rect 166 2116 220 2250
rect 220 2116 358 2250
rect 358 2116 412 2250
rect 412 2116 420 2250
rect 1150 2116 1180 2250
rect 1180 2116 1570 2250
rect 0 1882 420 2116
rect 1150 1882 1570 2116
rect 0 1750 166 1882
rect 166 1750 220 1882
rect 220 1750 358 1882
rect 358 1750 412 1882
rect 412 1750 420 1882
rect 1150 1750 1180 1882
rect 1180 1750 1570 1882
rect 520 1480 646 1610
rect 646 1480 700 1610
rect 700 1480 838 1610
rect 838 1480 892 1610
rect 892 1480 1030 1610
rect 1030 1480 1040 1610
rect 520 1450 1040 1480
rect 520 1246 1040 1270
rect 520 1110 646 1246
rect 646 1110 700 1246
rect 700 1110 838 1246
rect 838 1110 892 1246
rect 892 1110 1030 1246
rect 1030 1110 1040 1246
rect 0 844 166 980
rect 166 844 220 980
rect 220 844 358 980
rect 358 844 412 980
rect 412 844 420 980
rect 1150 844 1180 980
rect 1180 844 1570 980
rect 0 740 420 844
rect 1150 740 1570 844
rect 520 610 1040 640
rect 520 480 550 610
rect 550 480 604 610
rect 604 480 742 610
rect 742 480 796 610
rect 796 480 934 610
rect 934 480 988 610
rect 988 480 1040 610
rect 0 208 70 340
rect 70 208 124 340
rect 124 208 262 340
rect 262 208 316 340
rect 316 208 420 340
rect 1150 208 1222 340
rect 1222 208 1276 340
rect 1276 208 1570 340
rect 0 100 420 208
rect 1150 100 1570 208
<< metal3 >>
rect -10 4160 430 4165
rect -10 3840 0 4160
rect 420 3840 430 4160
rect -10 3835 430 3840
rect 1140 4160 1580 4165
rect 1140 3840 1150 4160
rect 1570 3840 1580 4160
rect 1140 3835 1580 3840
rect 0 3475 420 3835
rect 520 3715 1040 3720
rect 510 3710 1050 3715
rect 510 3550 520 3710
rect 1040 3550 1050 3710
rect 510 3545 1050 3550
rect -10 3470 430 3475
rect -10 3210 0 3470
rect 420 3210 430 3470
rect -10 3205 430 3210
rect 0 3200 420 3205
rect 520 3075 1040 3545
rect 1150 3475 1570 3835
rect 1140 3470 1580 3475
rect 1140 3210 1150 3470
rect 1570 3210 1580 3470
rect 1140 3205 1580 3210
rect 1150 3200 1570 3205
rect 510 3070 1050 3075
rect 510 2910 520 3070
rect 1040 2910 1050 3070
rect 510 2905 1050 2910
rect 520 2545 1040 2905
rect 510 2540 1050 2545
rect 510 2380 520 2540
rect 1040 2380 1050 2540
rect 510 2375 1050 2380
rect 0 2255 420 2260
rect -10 2250 430 2255
rect -10 1750 0 2250
rect 420 1750 430 2250
rect -10 1745 430 1750
rect 0 985 420 1745
rect 520 1615 1040 2375
rect 1150 2255 1570 2260
rect 1140 2250 1580 2255
rect 1140 1750 1150 2250
rect 1570 1750 1580 2250
rect 1140 1745 1580 1750
rect 510 1610 1050 1615
rect 510 1450 520 1610
rect 1040 1450 1050 1610
rect 510 1445 1050 1450
rect 520 1275 1040 1445
rect 510 1270 1050 1275
rect 510 1110 520 1270
rect 1040 1110 1050 1270
rect 510 1105 1050 1110
rect -10 980 430 985
rect -10 740 0 980
rect 420 740 430 980
rect -10 735 430 740
rect 0 345 420 735
rect 520 645 1040 1105
rect 1150 985 1570 1745
rect 1140 980 1580 985
rect 1140 740 1150 980
rect 1570 740 1580 980
rect 1140 735 1580 740
rect 510 640 1050 645
rect 510 480 520 640
rect 1040 480 1050 640
rect 510 475 1050 480
rect 520 470 1040 475
rect 1150 345 1570 735
rect -10 340 430 345
rect -10 100 0 340
rect 420 100 430 340
rect -10 95 430 100
rect 1140 340 1580 345
rect 1140 100 1150 340
rect 1570 100 1580 340
rect 1140 95 1580 100
rect 0 80 420 95
rect 1150 80 1570 95
use sky130_fd_pr__pfet_01v8_8DK6RJ  sky130_fd_pr__pfet_01v8_8DK6RJ_0
timestamp 1654768133
transform 1 0 673 0 1 1363
box -743 -1373 743 1373
use sky130_fd_pr__pfet_01v8_9Z5L4S  sky130_fd_pr__pfet_01v8_9Z5L4S_0
timestamp 1654768133
transform 1 0 805 0 -1 3457
box -875 -737 875 737
<< end >>
