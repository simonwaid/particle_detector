magic
tech sky130B
magscale 1 2
timestamp 1654002310
<< error_p >>
rect -317 272 -259 278
rect -125 272 -67 278
rect 67 272 125 278
rect 259 272 317 278
rect -317 238 -305 272
rect -125 238 -113 272
rect 67 238 79 272
rect 259 238 271 272
rect -317 232 -259 238
rect -125 232 -67 238
rect 67 232 125 238
rect 259 232 317 238
rect -413 -238 -355 -232
rect -221 -238 -163 -232
rect -29 -238 29 -232
rect 163 -238 221 -232
rect 355 -238 413 -232
rect -413 -272 -401 -238
rect -221 -272 -209 -238
rect -29 -272 -17 -238
rect 163 -272 175 -238
rect 355 -272 367 -238
rect -413 -278 -355 -272
rect -221 -278 -163 -272
rect -29 -278 29 -272
rect 163 -278 221 -272
rect 355 -278 413 -272
<< pwell >>
rect -599 -410 599 410
<< nmoslvt >>
rect -399 -200 -369 200
rect -303 -200 -273 200
rect -207 -200 -177 200
rect -111 -200 -81 200
rect -15 -200 15 200
rect 81 -200 111 200
rect 177 -200 207 200
rect 273 -200 303 200
rect 369 -200 399 200
<< ndiff >>
rect -461 188 -399 200
rect -461 -188 -449 188
rect -415 -188 -399 188
rect -461 -200 -399 -188
rect -369 188 -303 200
rect -369 -188 -353 188
rect -319 -188 -303 188
rect -369 -200 -303 -188
rect -273 188 -207 200
rect -273 -188 -257 188
rect -223 -188 -207 188
rect -273 -200 -207 -188
rect -177 188 -111 200
rect -177 -188 -161 188
rect -127 -188 -111 188
rect -177 -200 -111 -188
rect -81 188 -15 200
rect -81 -188 -65 188
rect -31 -188 -15 188
rect -81 -200 -15 -188
rect 15 188 81 200
rect 15 -188 31 188
rect 65 -188 81 188
rect 15 -200 81 -188
rect 111 188 177 200
rect 111 -188 127 188
rect 161 -188 177 188
rect 111 -200 177 -188
rect 207 188 273 200
rect 207 -188 223 188
rect 257 -188 273 188
rect 207 -200 273 -188
rect 303 188 369 200
rect 303 -188 319 188
rect 353 -188 369 188
rect 303 -200 369 -188
rect 399 188 461 200
rect 399 -188 415 188
rect 449 -188 461 188
rect 399 -200 461 -188
<< ndiffc >>
rect -449 -188 -415 188
rect -353 -188 -319 188
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
rect 319 -188 353 188
rect 415 -188 449 188
<< psubdiff >>
rect -563 340 -467 374
rect 467 340 563 374
rect -563 278 -529 340
rect 529 278 563 340
rect -563 -340 -529 -278
rect 529 -340 563 -278
rect -563 -374 -467 -340
rect 467 -374 563 -340
<< psubdiffcont >>
rect -467 340 467 374
rect -563 -278 -529 278
rect 529 -278 563 278
rect -467 -374 467 -340
<< poly >>
rect -321 272 -255 288
rect -321 238 -305 272
rect -271 238 -255 272
rect -399 200 -369 226
rect -321 222 -255 238
rect -129 272 -63 288
rect -129 238 -113 272
rect -79 238 -63 272
rect -303 200 -273 222
rect -207 200 -177 226
rect -129 222 -63 238
rect 63 272 129 288
rect 63 238 79 272
rect 113 238 129 272
rect -111 200 -81 222
rect -15 200 15 226
rect 63 222 129 238
rect 255 272 321 288
rect 255 238 271 272
rect 305 238 321 272
rect 81 200 111 222
rect 177 200 207 226
rect 255 222 321 238
rect 273 200 303 222
rect 369 200 399 226
rect -399 -222 -369 -200
rect -417 -238 -351 -222
rect -303 -226 -273 -200
rect -207 -222 -177 -200
rect -417 -272 -401 -238
rect -367 -272 -351 -238
rect -417 -288 -351 -272
rect -225 -238 -159 -222
rect -111 -226 -81 -200
rect -15 -222 15 -200
rect -225 -272 -209 -238
rect -175 -272 -159 -238
rect -225 -288 -159 -272
rect -33 -238 33 -222
rect 81 -226 111 -200
rect 177 -222 207 -200
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
rect 159 -238 225 -222
rect 273 -226 303 -200
rect 369 -222 399 -200
rect 159 -272 175 -238
rect 209 -272 225 -238
rect 159 -288 225 -272
rect 351 -238 417 -222
rect 351 -272 367 -238
rect 401 -272 417 -238
rect 351 -288 417 -272
<< polycont >>
rect -305 238 -271 272
rect -113 238 -79 272
rect 79 238 113 272
rect 271 238 305 272
rect -401 -272 -367 -238
rect -209 -272 -175 -238
rect -17 -272 17 -238
rect 175 -272 209 -238
rect 367 -272 401 -238
<< locali >>
rect -563 340 -467 374
rect 467 340 563 374
rect -563 278 -529 340
rect 529 278 563 340
rect -321 238 -305 272
rect -271 238 -255 272
rect -129 238 -113 272
rect -79 238 -63 272
rect 63 238 79 272
rect 113 238 129 272
rect 255 238 271 272
rect 305 238 321 272
rect -449 188 -415 204
rect -449 -204 -415 -188
rect -353 188 -319 204
rect -353 -204 -319 -188
rect -257 188 -223 204
rect -257 -204 -223 -188
rect -161 188 -127 204
rect -161 -204 -127 -188
rect -65 188 -31 204
rect -65 -204 -31 -188
rect 31 188 65 204
rect 31 -204 65 -188
rect 127 188 161 204
rect 127 -204 161 -188
rect 223 188 257 204
rect 223 -204 257 -188
rect 319 188 353 204
rect 319 -204 353 -188
rect 415 188 449 204
rect 415 -204 449 -188
rect -417 -272 -401 -238
rect -367 -272 -351 -238
rect -225 -272 -209 -238
rect -175 -272 -159 -238
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 159 -272 175 -238
rect 209 -272 225 -238
rect 351 -272 367 -238
rect 401 -272 417 -238
rect -563 -340 -529 -278
rect 529 -340 563 -278
rect -563 -374 -467 -340
rect 467 -374 563 -340
<< viali >>
rect -305 238 -271 272
rect -113 238 -79 272
rect 79 238 113 272
rect 271 238 305 272
rect -449 -188 -415 188
rect -353 -188 -319 188
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
rect 319 -188 353 188
rect 415 -188 449 188
rect -401 -272 -367 -238
rect -209 -272 -175 -238
rect -17 -272 17 -238
rect 175 -272 209 -238
rect 367 -272 401 -238
<< metal1 >>
rect -317 272 -259 278
rect -317 238 -305 272
rect -271 238 -259 272
rect -317 232 -259 238
rect -125 272 -67 278
rect -125 238 -113 272
rect -79 238 -67 272
rect -125 232 -67 238
rect 67 272 125 278
rect 67 238 79 272
rect 113 238 125 272
rect 67 232 125 238
rect 259 272 317 278
rect 259 238 271 272
rect 305 238 317 272
rect 259 232 317 238
rect -455 188 -409 200
rect -455 -188 -449 188
rect -415 -188 -409 188
rect -455 -200 -409 -188
rect -359 188 -313 200
rect -359 -188 -353 188
rect -319 -188 -313 188
rect -359 -200 -313 -188
rect -263 188 -217 200
rect -263 -188 -257 188
rect -223 -188 -217 188
rect -263 -200 -217 -188
rect -167 188 -121 200
rect -167 -188 -161 188
rect -127 -188 -121 188
rect -167 -200 -121 -188
rect -71 188 -25 200
rect -71 -188 -65 188
rect -31 -188 -25 188
rect -71 -200 -25 -188
rect 25 188 71 200
rect 25 -188 31 188
rect 65 -188 71 188
rect 25 -200 71 -188
rect 121 188 167 200
rect 121 -188 127 188
rect 161 -188 167 188
rect 121 -200 167 -188
rect 217 188 263 200
rect 217 -188 223 188
rect 257 -188 263 188
rect 217 -200 263 -188
rect 313 188 359 200
rect 313 -188 319 188
rect 353 -188 359 188
rect 313 -200 359 -188
rect 409 188 455 200
rect 409 -188 415 188
rect 449 -188 455 188
rect 409 -200 455 -188
rect -413 -238 -355 -232
rect -413 -272 -401 -238
rect -367 -272 -355 -238
rect -413 -278 -355 -272
rect -221 -238 -163 -232
rect -221 -272 -209 -238
rect -175 -272 -163 -238
rect -221 -278 -163 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 163 -238 221 -232
rect 163 -272 175 -238
rect 209 -272 221 -238
rect 163 -278 221 -272
rect 355 -238 413 -232
rect 355 -272 367 -238
rect 401 -272 413 -238
rect 355 -278 413 -272
<< properties >>
string FIXED_BBOX -546 -357 546 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 1 nf 9 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
