magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< metal1 >>
rect 620 110 880 160
rect 900 120 1210 180
rect 2000 120 2310 180
rect 3050 120 3360 180
rect 4110 120 4420 180
rect 5250 120 5560 180
rect 6330 120 6640 180
rect 7420 120 7730 180
rect 8510 120 8820 180
rect 620 30 630 110
rect 870 30 880 110
<< via1 >>
rect 630 30 870 110
<< metal2 >>
rect 290 2240 610 2250
rect 290 1950 610 1960
rect 1380 2240 1700 2250
rect 1380 1950 1700 1960
rect 2460 2240 2780 2250
rect 2460 1950 2780 1960
rect 3550 2240 3870 2250
rect 3550 1950 3870 1960
rect 4640 2240 4960 2250
rect 4640 1950 4960 1960
rect 5730 2240 6050 2250
rect 5730 1950 6050 1960
rect 6820 2240 7140 2250
rect 6820 1950 7140 1960
rect 7910 2240 8230 2250
rect 7910 1950 8230 1960
rect 9000 2240 9320 2250
rect 9000 1950 9320 1960
rect 630 110 870 120
rect 630 20 870 30
<< via2 >>
rect 290 1960 610 2240
rect 1380 1960 1700 2240
rect 2460 1960 2780 2240
rect 3550 1960 3870 2240
rect 4640 1960 4960 2240
rect 5730 1960 6050 2240
rect 6820 1960 7140 2240
rect 7910 1960 8230 2240
rect 9000 1960 9320 2240
rect 630 30 870 110
<< metal3 >>
rect 280 2240 620 2245
rect 280 1960 290 2240
rect 610 1960 620 2240
rect 280 1955 620 1960
rect 1370 2240 1710 2245
rect 1370 1960 1380 2240
rect 1700 1960 1710 2240
rect 1370 1955 1710 1960
rect 2450 2240 2790 2245
rect 2450 1960 2460 2240
rect 2780 1960 2790 2240
rect 2450 1955 2790 1960
rect 3540 2240 3880 2245
rect 3540 1960 3550 2240
rect 3870 1960 3880 2240
rect 3540 1955 3880 1960
rect 4630 2240 4970 2245
rect 4630 1960 4640 2240
rect 4960 1960 4970 2240
rect 4630 1955 4970 1960
rect 5720 2240 6060 2245
rect 5720 1960 5730 2240
rect 6050 1960 6060 2240
rect 5720 1955 6060 1960
rect 6810 2240 7150 2245
rect 6810 1960 6820 2240
rect 7140 1960 7150 2240
rect 6810 1955 7150 1960
rect 7900 2240 8240 2245
rect 7900 1960 7910 2240
rect 8230 1960 8240 2240
rect 7900 1955 8240 1960
rect 8990 2240 9330 2245
rect 8990 1960 9000 2240
rect 9320 1960 9330 2240
rect 8990 1955 9330 1960
rect 630 115 870 620
rect 620 110 880 115
rect 620 30 630 110
rect 870 30 880 110
rect 1720 60 1960 620
rect 2810 60 3050 620
rect 3900 60 4140 620
rect 4990 60 5230 620
rect 6080 60 6320 620
rect 7170 60 7410 620
rect 8260 60 8500 620
rect 9350 60 9590 620
rect 620 25 880 30
<< via3 >>
rect 290 1960 610 2240
rect 1380 1960 1700 2240
rect 2460 1960 2780 2240
rect 3550 1960 3870 2240
rect 4640 1960 4960 2240
rect 5730 1960 6050 2240
rect 6820 1960 7140 2240
rect 7910 1960 8230 2240
rect 9000 1960 9320 2240
<< metal4 >>
rect 289 2240 611 2241
rect 289 1960 290 2240
rect 610 1960 611 2240
rect 289 1959 611 1960
rect 1379 2240 1701 2241
rect 1379 1960 1380 2240
rect 1700 1960 1701 2240
rect 1379 1959 1701 1960
rect 2459 2240 2781 2241
rect 2459 1960 2460 2240
rect 2780 1960 2781 2240
rect 2459 1959 2781 1960
rect 3549 2240 3871 2241
rect 3549 1960 3550 2240
rect 3870 1960 3871 2240
rect 3549 1959 3871 1960
rect 4639 2240 4961 2241
rect 4639 1960 4640 2240
rect 4960 1960 4961 2240
rect 4639 1959 4961 1960
rect 5729 2240 6051 2241
rect 5729 1960 5730 2240
rect 6050 1960 6051 2240
rect 5729 1959 6051 1960
rect 6819 2240 7141 2241
rect 6819 1960 6820 2240
rect 7140 1960 7141 2240
rect 6819 1959 7141 1960
rect 7909 2240 8231 2241
rect 7909 1960 7910 2240
rect 8230 1960 8231 2240
rect 7909 1959 8231 1960
rect 8999 2240 9321 2241
rect 8999 1960 9000 2240
rect 9320 1960 9321 2240
rect 8999 1959 9321 1960
<< via4 >>
rect 290 1960 610 2240
rect 1380 1960 1700 2240
rect 2460 1960 2780 2240
rect 3550 1960 3870 2240
rect 4640 1960 4960 2240
rect 5730 1960 6050 2240
rect 6820 1960 7140 2240
rect 7910 1960 8230 2240
rect 9000 1960 9320 2240
<< metal5 >>
rect 0 2240 9830 2300
rect 0 1960 290 2240
rect 610 1960 1380 2240
rect 1700 1960 2460 2240
rect 2780 1960 3550 2240
rect 3870 1960 4640 2240
rect 4960 1960 5730 2240
rect 6050 1960 6820 2240
rect 7140 1960 7910 2240
rect 8230 1960 9000 2240
rect 9320 1960 9830 2240
rect 0 1940 9830 1960
rect 266 1936 634 1940
rect 1356 1936 1724 1940
rect 2436 1936 2804 1940
rect 3526 1936 3894 1940
rect 4616 1936 4984 1940
rect 5706 1936 6074 1940
rect 6796 1936 7164 1940
rect 7886 1936 8254 1940
rect 8976 1936 9344 1940
use bias_curm_p  bias_curm_p_0
timestamp 1654760956
transform 1 0 10 0 1 910
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_1
timestamp 1654760956
transform 1 0 1100 0 1 910
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_2
timestamp 1654760956
transform 1 0 2190 0 1 910
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_3
timestamp 1654760956
transform 1 0 3280 0 1 910
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_4
timestamp 1654760956
transform 1 0 6550 0 1 910
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_5
timestamp 1654760956
transform 1 0 5460 0 1 910
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_6
timestamp 1654760956
transform 1 0 4370 0 1 910
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_7
timestamp 1654760956
transform 1 0 8730 0 1 910
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_8
timestamp 1654760956
transform 1 0 7640 0 1 910
box -10 -910 1100 1390
<< labels >>
rlabel metal3 680 60 790 150 1 I_in
rlabel space 1750 50 1860 140 1 I_out1
rlabel metal3 2850 60 2960 150 1 I_out2
rlabel metal3 3940 70 4050 160 1 I_out3
rlabel metal3 5030 70 5140 160 1 I_out4
rlabel metal3 6130 70 6240 160 1 I_out5
rlabel metal3 7200 70 7310 160 1 I_out6
rlabel metal3 8290 70 8400 160 1 I_out7
rlabel metal3 9400 70 9510 160 1 I_out8
<< end >>
