magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< error_p >>
rect -678 599 -620 605
rect -560 599 -502 605
rect -442 599 -384 605
rect -324 599 -266 605
rect -206 599 -148 605
rect -88 599 -30 605
rect 30 599 88 605
rect 148 599 206 605
rect 266 599 324 605
rect 384 599 442 605
rect 502 599 560 605
rect 620 599 678 605
rect -678 565 -666 599
rect -560 565 -548 599
rect -442 565 -430 599
rect -324 565 -312 599
rect -206 565 -194 599
rect -88 565 -76 599
rect 30 565 42 599
rect 148 565 160 599
rect 266 565 278 599
rect 384 565 396 599
rect 502 565 514 599
rect 620 565 632 599
rect -678 559 -620 565
rect -560 559 -502 565
rect -442 559 -384 565
rect -324 559 -266 565
rect -206 559 -148 565
rect -88 559 -30 565
rect 30 559 88 565
rect 148 559 206 565
rect 266 559 324 565
rect 384 559 442 565
rect 502 559 560 565
rect 620 559 678 565
rect -678 71 -620 77
rect -560 71 -502 77
rect -442 71 -384 77
rect -324 71 -266 77
rect -206 71 -148 77
rect -88 71 -30 77
rect 30 71 88 77
rect 148 71 206 77
rect 266 71 324 77
rect 384 71 442 77
rect 502 71 560 77
rect 620 71 678 77
rect -678 37 -666 71
rect -560 37 -548 71
rect -442 37 -430 71
rect -324 37 -312 71
rect -206 37 -194 71
rect -88 37 -76 71
rect 30 37 42 71
rect 148 37 160 71
rect 266 37 278 71
rect 384 37 396 71
rect 502 37 514 71
rect 620 37 632 71
rect -678 31 -620 37
rect -560 31 -502 37
rect -442 31 -384 37
rect -324 31 -266 37
rect -206 31 -148 37
rect -88 31 -30 37
rect 30 31 88 37
rect 148 31 206 37
rect 266 31 324 37
rect 384 31 442 37
rect 502 31 560 37
rect 620 31 678 37
rect -678 -37 -620 -31
rect -560 -37 -502 -31
rect -442 -37 -384 -31
rect -324 -37 -266 -31
rect -206 -37 -148 -31
rect -88 -37 -30 -31
rect 30 -37 88 -31
rect 148 -37 206 -31
rect 266 -37 324 -31
rect 384 -37 442 -31
rect 502 -37 560 -31
rect 620 -37 678 -31
rect -678 -71 -666 -37
rect -560 -71 -548 -37
rect -442 -71 -430 -37
rect -324 -71 -312 -37
rect -206 -71 -194 -37
rect -88 -71 -76 -37
rect 30 -71 42 -37
rect 148 -71 160 -37
rect 266 -71 278 -37
rect 384 -71 396 -37
rect 502 -71 514 -37
rect 620 -71 632 -37
rect -678 -77 -620 -71
rect -560 -77 -502 -71
rect -442 -77 -384 -71
rect -324 -77 -266 -71
rect -206 -77 -148 -71
rect -88 -77 -30 -71
rect 30 -77 88 -71
rect 148 -77 206 -71
rect 266 -77 324 -71
rect 384 -77 442 -71
rect 502 -77 560 -71
rect 620 -77 678 -71
rect -678 -565 -620 -559
rect -560 -565 -502 -559
rect -442 -565 -384 -559
rect -324 -565 -266 -559
rect -206 -565 -148 -559
rect -88 -565 -30 -559
rect 30 -565 88 -559
rect 148 -565 206 -559
rect 266 -565 324 -559
rect 384 -565 442 -559
rect 502 -565 560 -559
rect 620 -565 678 -559
rect -678 -599 -666 -565
rect -560 -599 -548 -565
rect -442 -599 -430 -565
rect -324 -599 -312 -565
rect -206 -599 -194 -565
rect -88 -599 -76 -565
rect 30 -599 42 -565
rect 148 -599 160 -565
rect 266 -599 278 -565
rect 384 -599 396 -565
rect 502 -599 514 -565
rect 620 -599 632 -565
rect -678 -605 -620 -599
rect -560 -605 -502 -599
rect -442 -605 -384 -599
rect -324 -605 -266 -599
rect -206 -605 -148 -599
rect -88 -605 -30 -599
rect 30 -605 88 -599
rect 148 -605 206 -599
rect 266 -605 324 -599
rect 384 -605 442 -599
rect 502 -605 560 -599
rect 620 -605 678 -599
<< nwell >>
rect -875 -737 875 737
<< pmos >>
rect -679 118 -619 518
rect -561 118 -501 518
rect -443 118 -383 518
rect -325 118 -265 518
rect -207 118 -147 518
rect -89 118 -29 518
rect 29 118 89 518
rect 147 118 207 518
rect 265 118 325 518
rect 383 118 443 518
rect 501 118 561 518
rect 619 118 679 518
rect -679 -518 -619 -118
rect -561 -518 -501 -118
rect -443 -518 -383 -118
rect -325 -518 -265 -118
rect -207 -518 -147 -118
rect -89 -518 -29 -118
rect 29 -518 89 -118
rect 147 -518 207 -118
rect 265 -518 325 -118
rect 383 -518 443 -118
rect 501 -518 561 -118
rect 619 -518 679 -118
<< pdiff >>
rect -737 506 -679 518
rect -737 130 -725 506
rect -691 130 -679 506
rect -737 118 -679 130
rect -619 506 -561 518
rect -619 130 -607 506
rect -573 130 -561 506
rect -619 118 -561 130
rect -501 506 -443 518
rect -501 130 -489 506
rect -455 130 -443 506
rect -501 118 -443 130
rect -383 506 -325 518
rect -383 130 -371 506
rect -337 130 -325 506
rect -383 118 -325 130
rect -265 506 -207 518
rect -265 130 -253 506
rect -219 130 -207 506
rect -265 118 -207 130
rect -147 506 -89 518
rect -147 130 -135 506
rect -101 130 -89 506
rect -147 118 -89 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 89 506 147 518
rect 89 130 101 506
rect 135 130 147 506
rect 89 118 147 130
rect 207 506 265 518
rect 207 130 219 506
rect 253 130 265 506
rect 207 118 265 130
rect 325 506 383 518
rect 325 130 337 506
rect 371 130 383 506
rect 325 118 383 130
rect 443 506 501 518
rect 443 130 455 506
rect 489 130 501 506
rect 443 118 501 130
rect 561 506 619 518
rect 561 130 573 506
rect 607 130 619 506
rect 561 118 619 130
rect 679 506 737 518
rect 679 130 691 506
rect 725 130 737 506
rect 679 118 737 130
rect -737 -130 -679 -118
rect -737 -506 -725 -130
rect -691 -506 -679 -130
rect -737 -518 -679 -506
rect -619 -130 -561 -118
rect -619 -506 -607 -130
rect -573 -506 -561 -130
rect -619 -518 -561 -506
rect -501 -130 -443 -118
rect -501 -506 -489 -130
rect -455 -506 -443 -130
rect -501 -518 -443 -506
rect -383 -130 -325 -118
rect -383 -506 -371 -130
rect -337 -506 -325 -130
rect -383 -518 -325 -506
rect -265 -130 -207 -118
rect -265 -506 -253 -130
rect -219 -506 -207 -130
rect -265 -518 -207 -506
rect -147 -130 -89 -118
rect -147 -506 -135 -130
rect -101 -506 -89 -130
rect -147 -518 -89 -506
rect -29 -130 29 -118
rect -29 -506 -17 -130
rect 17 -506 29 -130
rect -29 -518 29 -506
rect 89 -130 147 -118
rect 89 -506 101 -130
rect 135 -506 147 -130
rect 89 -518 147 -506
rect 207 -130 265 -118
rect 207 -506 219 -130
rect 253 -506 265 -130
rect 207 -518 265 -506
rect 325 -130 383 -118
rect 325 -506 337 -130
rect 371 -506 383 -130
rect 325 -518 383 -506
rect 443 -130 501 -118
rect 443 -506 455 -130
rect 489 -506 501 -130
rect 443 -518 501 -506
rect 561 -130 619 -118
rect 561 -506 573 -130
rect 607 -506 619 -130
rect 561 -518 619 -506
rect 679 -130 737 -118
rect 679 -506 691 -130
rect 725 -506 737 -130
rect 679 -518 737 -506
<< pdiffc >>
rect -725 130 -691 506
rect -607 130 -573 506
rect -489 130 -455 506
rect -371 130 -337 506
rect -253 130 -219 506
rect -135 130 -101 506
rect -17 130 17 506
rect 101 130 135 506
rect 219 130 253 506
rect 337 130 371 506
rect 455 130 489 506
rect 573 130 607 506
rect 691 130 725 506
rect -725 -506 -691 -130
rect -607 -506 -573 -130
rect -489 -506 -455 -130
rect -371 -506 -337 -130
rect -253 -506 -219 -130
rect -135 -506 -101 -130
rect -17 -506 17 -130
rect 101 -506 135 -130
rect 219 -506 253 -130
rect 337 -506 371 -130
rect 455 -506 489 -130
rect 573 -506 607 -130
rect 691 -506 725 -130
<< nsubdiff >>
rect -839 667 -743 701
rect 743 667 839 701
rect -839 605 -805 667
rect 805 605 839 667
rect -839 -667 -805 -605
rect 805 -667 839 -605
rect -839 -701 -743 -667
rect 743 -701 839 -667
<< nsubdiffcont >>
rect -743 667 743 701
rect -839 -605 -805 605
rect 805 -605 839 605
rect -743 -701 743 -667
<< poly >>
rect -682 599 -616 615
rect -682 565 -666 599
rect -632 565 -616 599
rect -682 549 -616 565
rect -564 599 -498 615
rect -564 565 -548 599
rect -514 565 -498 599
rect -564 549 -498 565
rect -446 599 -380 615
rect -446 565 -430 599
rect -396 565 -380 599
rect -446 549 -380 565
rect -328 599 -262 615
rect -328 565 -312 599
rect -278 565 -262 599
rect -328 549 -262 565
rect -210 599 -144 615
rect -210 565 -194 599
rect -160 565 -144 599
rect -210 549 -144 565
rect -92 599 -26 615
rect -92 565 -76 599
rect -42 565 -26 599
rect -92 549 -26 565
rect 26 599 92 615
rect 26 565 42 599
rect 76 565 92 599
rect 26 549 92 565
rect 144 599 210 615
rect 144 565 160 599
rect 194 565 210 599
rect 144 549 210 565
rect 262 599 328 615
rect 262 565 278 599
rect 312 565 328 599
rect 262 549 328 565
rect 380 599 446 615
rect 380 565 396 599
rect 430 565 446 599
rect 380 549 446 565
rect 498 599 564 615
rect 498 565 514 599
rect 548 565 564 599
rect 498 549 564 565
rect 616 599 682 615
rect 616 565 632 599
rect 666 565 682 599
rect 616 549 682 565
rect -679 518 -619 549
rect -561 518 -501 549
rect -443 518 -383 549
rect -325 518 -265 549
rect -207 518 -147 549
rect -89 518 -29 549
rect 29 518 89 549
rect 147 518 207 549
rect 265 518 325 549
rect 383 518 443 549
rect 501 518 561 549
rect 619 518 679 549
rect -679 87 -619 118
rect -561 87 -501 118
rect -443 87 -383 118
rect -325 87 -265 118
rect -207 87 -147 118
rect -89 87 -29 118
rect 29 87 89 118
rect 147 87 207 118
rect 265 87 325 118
rect 383 87 443 118
rect 501 87 561 118
rect 619 87 679 118
rect -682 71 -616 87
rect -682 37 -666 71
rect -632 37 -616 71
rect -682 21 -616 37
rect -564 71 -498 87
rect -564 37 -548 71
rect -514 37 -498 71
rect -564 21 -498 37
rect -446 71 -380 87
rect -446 37 -430 71
rect -396 37 -380 71
rect -446 21 -380 37
rect -328 71 -262 87
rect -328 37 -312 71
rect -278 37 -262 71
rect -328 21 -262 37
rect -210 71 -144 87
rect -210 37 -194 71
rect -160 37 -144 71
rect -210 21 -144 37
rect -92 71 -26 87
rect -92 37 -76 71
rect -42 37 -26 71
rect -92 21 -26 37
rect 26 71 92 87
rect 26 37 42 71
rect 76 37 92 71
rect 26 21 92 37
rect 144 71 210 87
rect 144 37 160 71
rect 194 37 210 71
rect 144 21 210 37
rect 262 71 328 87
rect 262 37 278 71
rect 312 37 328 71
rect 262 21 328 37
rect 380 71 446 87
rect 380 37 396 71
rect 430 37 446 71
rect 380 21 446 37
rect 498 71 564 87
rect 498 37 514 71
rect 548 37 564 71
rect 498 21 564 37
rect 616 71 682 87
rect 616 37 632 71
rect 666 37 682 71
rect 616 21 682 37
rect -682 -37 -616 -21
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -682 -87 -616 -71
rect -564 -37 -498 -21
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -564 -87 -498 -71
rect -446 -37 -380 -21
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -446 -87 -380 -71
rect -328 -37 -262 -21
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -328 -87 -262 -71
rect -210 -37 -144 -21
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -210 -87 -144 -71
rect -92 -37 -26 -21
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect -92 -87 -26 -71
rect 26 -37 92 -21
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 26 -87 92 -71
rect 144 -37 210 -21
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 144 -87 210 -71
rect 262 -37 328 -21
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 262 -87 328 -71
rect 380 -37 446 -21
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 380 -87 446 -71
rect 498 -37 564 -21
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 498 -87 564 -71
rect 616 -37 682 -21
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 616 -87 682 -71
rect -679 -118 -619 -87
rect -561 -118 -501 -87
rect -443 -118 -383 -87
rect -325 -118 -265 -87
rect -207 -118 -147 -87
rect -89 -118 -29 -87
rect 29 -118 89 -87
rect 147 -118 207 -87
rect 265 -118 325 -87
rect 383 -118 443 -87
rect 501 -118 561 -87
rect 619 -118 679 -87
rect -679 -549 -619 -518
rect -561 -549 -501 -518
rect -443 -549 -383 -518
rect -325 -549 -265 -518
rect -207 -549 -147 -518
rect -89 -549 -29 -518
rect 29 -549 89 -518
rect 147 -549 207 -518
rect 265 -549 325 -518
rect 383 -549 443 -518
rect 501 -549 561 -518
rect 619 -549 679 -518
rect -682 -565 -616 -549
rect -682 -599 -666 -565
rect -632 -599 -616 -565
rect -682 -615 -616 -599
rect -564 -565 -498 -549
rect -564 -599 -548 -565
rect -514 -599 -498 -565
rect -564 -615 -498 -599
rect -446 -565 -380 -549
rect -446 -599 -430 -565
rect -396 -599 -380 -565
rect -446 -615 -380 -599
rect -328 -565 -262 -549
rect -328 -599 -312 -565
rect -278 -599 -262 -565
rect -328 -615 -262 -599
rect -210 -565 -144 -549
rect -210 -599 -194 -565
rect -160 -599 -144 -565
rect -210 -615 -144 -599
rect -92 -565 -26 -549
rect -92 -599 -76 -565
rect -42 -599 -26 -565
rect -92 -615 -26 -599
rect 26 -565 92 -549
rect 26 -599 42 -565
rect 76 -599 92 -565
rect 26 -615 92 -599
rect 144 -565 210 -549
rect 144 -599 160 -565
rect 194 -599 210 -565
rect 144 -615 210 -599
rect 262 -565 328 -549
rect 262 -599 278 -565
rect 312 -599 328 -565
rect 262 -615 328 -599
rect 380 -565 446 -549
rect 380 -599 396 -565
rect 430 -599 446 -565
rect 380 -615 446 -599
rect 498 -565 564 -549
rect 498 -599 514 -565
rect 548 -599 564 -565
rect 498 -615 564 -599
rect 616 -565 682 -549
rect 616 -599 632 -565
rect 666 -599 682 -565
rect 616 -615 682 -599
<< polycont >>
rect -666 565 -632 599
rect -548 565 -514 599
rect -430 565 -396 599
rect -312 565 -278 599
rect -194 565 -160 599
rect -76 565 -42 599
rect 42 565 76 599
rect 160 565 194 599
rect 278 565 312 599
rect 396 565 430 599
rect 514 565 548 599
rect 632 565 666 599
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect -666 -599 -632 -565
rect -548 -599 -514 -565
rect -430 -599 -396 -565
rect -312 -599 -278 -565
rect -194 -599 -160 -565
rect -76 -599 -42 -565
rect 42 -599 76 -565
rect 160 -599 194 -565
rect 278 -599 312 -565
rect 396 -599 430 -565
rect 514 -599 548 -565
rect 632 -599 666 -565
<< locali >>
rect -839 667 -743 701
rect 743 667 839 701
rect -839 605 -805 667
rect 805 605 839 667
rect -682 565 -666 599
rect -632 565 -616 599
rect -564 565 -548 599
rect -514 565 -498 599
rect -446 565 -430 599
rect -396 565 -380 599
rect -328 565 -312 599
rect -278 565 -262 599
rect -210 565 -194 599
rect -160 565 -144 599
rect -92 565 -76 599
rect -42 565 -26 599
rect 26 565 42 599
rect 76 565 92 599
rect 144 565 160 599
rect 194 565 210 599
rect 262 565 278 599
rect 312 565 328 599
rect 380 565 396 599
rect 430 565 446 599
rect 498 565 514 599
rect 548 565 564 599
rect 616 565 632 599
rect 666 565 682 599
rect -725 506 -691 522
rect -725 114 -691 130
rect -607 506 -573 522
rect -607 114 -573 130
rect -489 506 -455 522
rect -489 114 -455 130
rect -371 506 -337 522
rect -371 114 -337 130
rect -253 506 -219 522
rect -253 114 -219 130
rect -135 506 -101 522
rect -135 114 -101 130
rect -17 506 17 522
rect -17 114 17 130
rect 101 506 135 522
rect 101 114 135 130
rect 219 506 253 522
rect 219 114 253 130
rect 337 506 371 522
rect 337 114 371 130
rect 455 506 489 522
rect 455 114 489 130
rect 573 506 607 522
rect 573 114 607 130
rect 691 506 725 522
rect 691 114 725 130
rect -682 37 -666 71
rect -632 37 -616 71
rect -564 37 -548 71
rect -514 37 -498 71
rect -446 37 -430 71
rect -396 37 -380 71
rect -328 37 -312 71
rect -278 37 -262 71
rect -210 37 -194 71
rect -160 37 -144 71
rect -92 37 -76 71
rect -42 37 -26 71
rect 26 37 42 71
rect 76 37 92 71
rect 144 37 160 71
rect 194 37 210 71
rect 262 37 278 71
rect 312 37 328 71
rect 380 37 396 71
rect 430 37 446 71
rect 498 37 514 71
rect 548 37 564 71
rect 616 37 632 71
rect 666 37 682 71
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 616 -71 632 -37
rect 666 -71 682 -37
rect -725 -130 -691 -114
rect -725 -522 -691 -506
rect -607 -130 -573 -114
rect -607 -522 -573 -506
rect -489 -130 -455 -114
rect -489 -522 -455 -506
rect -371 -130 -337 -114
rect -371 -522 -337 -506
rect -253 -130 -219 -114
rect -253 -522 -219 -506
rect -135 -130 -101 -114
rect -135 -522 -101 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 101 -130 135 -114
rect 101 -522 135 -506
rect 219 -130 253 -114
rect 219 -522 253 -506
rect 337 -130 371 -114
rect 337 -522 371 -506
rect 455 -130 489 -114
rect 455 -522 489 -506
rect 573 -130 607 -114
rect 573 -522 607 -506
rect 691 -130 725 -114
rect 691 -522 725 -506
rect -682 -599 -666 -565
rect -632 -599 -616 -565
rect -564 -599 -548 -565
rect -514 -599 -498 -565
rect -446 -599 -430 -565
rect -396 -599 -380 -565
rect -328 -599 -312 -565
rect -278 -599 -262 -565
rect -210 -599 -194 -565
rect -160 -599 -144 -565
rect -92 -599 -76 -565
rect -42 -599 -26 -565
rect 26 -599 42 -565
rect 76 -599 92 -565
rect 144 -599 160 -565
rect 194 -599 210 -565
rect 262 -599 278 -565
rect 312 -599 328 -565
rect 380 -599 396 -565
rect 430 -599 446 -565
rect 498 -599 514 -565
rect 548 -599 564 -565
rect 616 -599 632 -565
rect 666 -599 682 -565
rect -839 -667 -805 -605
rect 805 -667 839 -605
rect -839 -701 -743 -667
rect 743 -701 839 -667
<< viali >>
rect -666 565 -632 599
rect -548 565 -514 599
rect -430 565 -396 599
rect -312 565 -278 599
rect -194 565 -160 599
rect -76 565 -42 599
rect 42 565 76 599
rect 160 565 194 599
rect 278 565 312 599
rect 396 565 430 599
rect 514 565 548 599
rect 632 565 666 599
rect -725 130 -691 506
rect -607 130 -573 506
rect -489 130 -455 506
rect -371 130 -337 506
rect -253 130 -219 506
rect -135 130 -101 506
rect -17 130 17 506
rect 101 130 135 506
rect 219 130 253 506
rect 337 130 371 506
rect 455 130 489 506
rect 573 130 607 506
rect 691 130 725 506
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect -725 -506 -691 -130
rect -607 -506 -573 -130
rect -489 -506 -455 -130
rect -371 -506 -337 -130
rect -253 -506 -219 -130
rect -135 -506 -101 -130
rect -17 -506 17 -130
rect 101 -506 135 -130
rect 219 -506 253 -130
rect 337 -506 371 -130
rect 455 -506 489 -130
rect 573 -506 607 -130
rect 691 -506 725 -130
rect -666 -599 -632 -565
rect -548 -599 -514 -565
rect -430 -599 -396 -565
rect -312 -599 -278 -565
rect -194 -599 -160 -565
rect -76 -599 -42 -565
rect 42 -599 76 -565
rect 160 -599 194 -565
rect 278 -599 312 -565
rect 396 -599 430 -565
rect 514 -599 548 -565
rect 632 -599 666 -565
<< metal1 >>
rect -678 599 -620 605
rect -678 565 -666 599
rect -632 565 -620 599
rect -678 559 -620 565
rect -560 599 -502 605
rect -560 565 -548 599
rect -514 565 -502 599
rect -560 559 -502 565
rect -442 599 -384 605
rect -442 565 -430 599
rect -396 565 -384 599
rect -442 559 -384 565
rect -324 599 -266 605
rect -324 565 -312 599
rect -278 565 -266 599
rect -324 559 -266 565
rect -206 599 -148 605
rect -206 565 -194 599
rect -160 565 -148 599
rect -206 559 -148 565
rect -88 599 -30 605
rect -88 565 -76 599
rect -42 565 -30 599
rect -88 559 -30 565
rect 30 599 88 605
rect 30 565 42 599
rect 76 565 88 599
rect 30 559 88 565
rect 148 599 206 605
rect 148 565 160 599
rect 194 565 206 599
rect 148 559 206 565
rect 266 599 324 605
rect 266 565 278 599
rect 312 565 324 599
rect 266 559 324 565
rect 384 599 442 605
rect 384 565 396 599
rect 430 565 442 599
rect 384 559 442 565
rect 502 599 560 605
rect 502 565 514 599
rect 548 565 560 599
rect 502 559 560 565
rect 620 599 678 605
rect 620 565 632 599
rect 666 565 678 599
rect 620 559 678 565
rect -731 506 -685 518
rect -731 130 -725 506
rect -691 130 -685 506
rect -731 118 -685 130
rect -613 506 -567 518
rect -613 130 -607 506
rect -573 130 -567 506
rect -613 118 -567 130
rect -495 506 -449 518
rect -495 130 -489 506
rect -455 130 -449 506
rect -495 118 -449 130
rect -377 506 -331 518
rect -377 130 -371 506
rect -337 130 -331 506
rect -377 118 -331 130
rect -259 506 -213 518
rect -259 130 -253 506
rect -219 130 -213 506
rect -259 118 -213 130
rect -141 506 -95 518
rect -141 130 -135 506
rect -101 130 -95 506
rect -141 118 -95 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 95 506 141 518
rect 95 130 101 506
rect 135 130 141 506
rect 95 118 141 130
rect 213 506 259 518
rect 213 130 219 506
rect 253 130 259 506
rect 213 118 259 130
rect 331 506 377 518
rect 331 130 337 506
rect 371 130 377 506
rect 331 118 377 130
rect 449 506 495 518
rect 449 130 455 506
rect 489 130 495 506
rect 449 118 495 130
rect 567 506 613 518
rect 567 130 573 506
rect 607 130 613 506
rect 567 118 613 130
rect 685 506 731 518
rect 685 130 691 506
rect 725 130 731 506
rect 685 118 731 130
rect -678 71 -620 77
rect -678 37 -666 71
rect -632 37 -620 71
rect -678 31 -620 37
rect -560 71 -502 77
rect -560 37 -548 71
rect -514 37 -502 71
rect -560 31 -502 37
rect -442 71 -384 77
rect -442 37 -430 71
rect -396 37 -384 71
rect -442 31 -384 37
rect -324 71 -266 77
rect -324 37 -312 71
rect -278 37 -266 71
rect -324 31 -266 37
rect -206 71 -148 77
rect -206 37 -194 71
rect -160 37 -148 71
rect -206 31 -148 37
rect -88 71 -30 77
rect -88 37 -76 71
rect -42 37 -30 71
rect -88 31 -30 37
rect 30 71 88 77
rect 30 37 42 71
rect 76 37 88 71
rect 30 31 88 37
rect 148 71 206 77
rect 148 37 160 71
rect 194 37 206 71
rect 148 31 206 37
rect 266 71 324 77
rect 266 37 278 71
rect 312 37 324 71
rect 266 31 324 37
rect 384 71 442 77
rect 384 37 396 71
rect 430 37 442 71
rect 384 31 442 37
rect 502 71 560 77
rect 502 37 514 71
rect 548 37 560 71
rect 502 31 560 37
rect 620 71 678 77
rect 620 37 632 71
rect 666 37 678 71
rect 620 31 678 37
rect -678 -37 -620 -31
rect -678 -71 -666 -37
rect -632 -71 -620 -37
rect -678 -77 -620 -71
rect -560 -37 -502 -31
rect -560 -71 -548 -37
rect -514 -71 -502 -37
rect -560 -77 -502 -71
rect -442 -37 -384 -31
rect -442 -71 -430 -37
rect -396 -71 -384 -37
rect -442 -77 -384 -71
rect -324 -37 -266 -31
rect -324 -71 -312 -37
rect -278 -71 -266 -37
rect -324 -77 -266 -71
rect -206 -37 -148 -31
rect -206 -71 -194 -37
rect -160 -71 -148 -37
rect -206 -77 -148 -71
rect -88 -37 -30 -31
rect -88 -71 -76 -37
rect -42 -71 -30 -37
rect -88 -77 -30 -71
rect 30 -37 88 -31
rect 30 -71 42 -37
rect 76 -71 88 -37
rect 30 -77 88 -71
rect 148 -37 206 -31
rect 148 -71 160 -37
rect 194 -71 206 -37
rect 148 -77 206 -71
rect 266 -37 324 -31
rect 266 -71 278 -37
rect 312 -71 324 -37
rect 266 -77 324 -71
rect 384 -37 442 -31
rect 384 -71 396 -37
rect 430 -71 442 -37
rect 384 -77 442 -71
rect 502 -37 560 -31
rect 502 -71 514 -37
rect 548 -71 560 -37
rect 502 -77 560 -71
rect 620 -37 678 -31
rect 620 -71 632 -37
rect 666 -71 678 -37
rect 620 -77 678 -71
rect -731 -130 -685 -118
rect -731 -506 -725 -130
rect -691 -506 -685 -130
rect -731 -518 -685 -506
rect -613 -130 -567 -118
rect -613 -506 -607 -130
rect -573 -506 -567 -130
rect -613 -518 -567 -506
rect -495 -130 -449 -118
rect -495 -506 -489 -130
rect -455 -506 -449 -130
rect -495 -518 -449 -506
rect -377 -130 -331 -118
rect -377 -506 -371 -130
rect -337 -506 -331 -130
rect -377 -518 -331 -506
rect -259 -130 -213 -118
rect -259 -506 -253 -130
rect -219 -506 -213 -130
rect -259 -518 -213 -506
rect -141 -130 -95 -118
rect -141 -506 -135 -130
rect -101 -506 -95 -130
rect -141 -518 -95 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 95 -130 141 -118
rect 95 -506 101 -130
rect 135 -506 141 -130
rect 95 -518 141 -506
rect 213 -130 259 -118
rect 213 -506 219 -130
rect 253 -506 259 -130
rect 213 -518 259 -506
rect 331 -130 377 -118
rect 331 -506 337 -130
rect 371 -506 377 -130
rect 331 -518 377 -506
rect 449 -130 495 -118
rect 449 -506 455 -130
rect 489 -506 495 -130
rect 449 -518 495 -506
rect 567 -130 613 -118
rect 567 -506 573 -130
rect 607 -506 613 -130
rect 567 -518 613 -506
rect 685 -130 731 -118
rect 685 -506 691 -130
rect 725 -506 731 -130
rect 685 -518 731 -506
rect -678 -565 -620 -559
rect -678 -599 -666 -565
rect -632 -599 -620 -565
rect -678 -605 -620 -599
rect -560 -565 -502 -559
rect -560 -599 -548 -565
rect -514 -599 -502 -565
rect -560 -605 -502 -599
rect -442 -565 -384 -559
rect -442 -599 -430 -565
rect -396 -599 -384 -565
rect -442 -605 -384 -599
rect -324 -565 -266 -559
rect -324 -599 -312 -565
rect -278 -599 -266 -565
rect -324 -605 -266 -599
rect -206 -565 -148 -559
rect -206 -599 -194 -565
rect -160 -599 -148 -565
rect -206 -605 -148 -599
rect -88 -565 -30 -559
rect -88 -599 -76 -565
rect -42 -599 -30 -565
rect -88 -605 -30 -599
rect 30 -565 88 -559
rect 30 -599 42 -565
rect 76 -599 88 -565
rect 30 -605 88 -599
rect 148 -565 206 -559
rect 148 -599 160 -565
rect 194 -599 206 -565
rect 148 -605 206 -599
rect 266 -565 324 -559
rect 266 -599 278 -565
rect 312 -599 324 -565
rect 266 -605 324 -599
rect 384 -565 442 -559
rect 384 -599 396 -565
rect 430 -599 442 -565
rect 384 -605 442 -599
rect 502 -565 560 -559
rect 502 -599 514 -565
rect 548 -599 560 -565
rect 502 -605 560 -599
rect 620 -565 678 -559
rect 620 -599 632 -565
rect 666 -599 678 -565
rect 620 -605 678 -599
<< properties >>
string FIXED_BBOX -822 -684 822 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.3 m 2 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
