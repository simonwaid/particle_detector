* SPICE3 file created from outd.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2 m4_n3351_n3100# c2_n3251_n3000#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WXTTNJ c1_n2050_n2000# m3_n2150_n2100#
X0 c1_n2050_n2000# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
.ends

.subckt sky130_fd_pr__res_high_po_5p73_PA2QZX a_n573_400# a_n573_n832# a_n703_n962#
X0 a_n573_n832# a_n573_400# a_n703_n962# sky130_fd_pr__res_high_po_5p73 l=4e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_324MKY a_n369_n509# a_n81_109# a_n129_531# a_303_n509#
+ a_351_n87# a_n33_n87# a_399_109# a_n129_n597# a_n513_n597# a_63_n597# a_n273_109#
+ a_n465_n509# a_n225_n87# a_447_531# a_15_109# a_n321_531# a_15_n509# a_n177_n509#
+ a_111_n509# a_n321_n597# a_207_109# a_n417_n87# a_n465_109# a_n273_n509# a_351_21#
+ a_n513_531# a_n33_21# a_n225_21# a_n177_109# a_447_n597# a_n557_n509# a_495_109#
+ a_399_n509# a_n81_n509# a_111_109# a_n557_109# a_n369_109# a_159_21# a_495_n509#
+ a_63_531# a_255_n597# a_n659_n683# a_159_n87# a_n417_21# a_303_109# a_255_531# a_207_n509#
X0 a_399_n509# a_351_n87# a_303_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n81_109# a_n129_531# a_n177_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_111_109# a_63_531# a_15_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_n465_n509# a_n513_n597# a_n557_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X4 a_n273_109# a_n321_531# a_n369_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_n177_109# a_n225_21# a_n273_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 a_n81_n509# a_n129_n597# a_n177_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_15_n509# a_n33_n87# a_n81_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X8 a_n369_n509# a_n417_n87# a_n465_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X9 a_303_n509# a_255_n597# a_207_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X10 a_n273_n509# a_n321_n597# a_n369_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_303_109# a_255_531# a_207_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_207_109# a_159_21# a_111_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 a_399_109# a_351_21# a_303_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X14 a_495_109# a_447_531# a_399_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X15 a_n177_n509# a_n225_n87# a_n273_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 a_207_n509# a_159_n87# a_111_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17 a_495_n509# a_447_n597# a_399_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X18 a_n465_109# a_n513_531# a_n557_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X19 a_n369_109# a_n417_21# a_n465_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 a_111_n509# a_63_n597# a_15_n509# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 a_15_109# a_n33_21# a_n81_109# a_n659_n683# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt outd_diffamp m1_610_8380# m1_226_8380# m1_802_8758# m1_418_8758# m1_2276_8758#
+ m1_2084_8380# m1_1700_8758# m1_1186_8380# m1_898_8998# m1_130_8998# m1_706_8140#
+ m1_1796_8998# m1_1090_8998# m1_2564_8140# m1_1604_8140# m1_610_8758# m1_226_8758#
+ m1_2084_8758# m1_1186_8758# m1_514_8140# m1_706_8998# m1_2564_8998# m1_2372_8140#
+ m1_1604_8998# m1_994_8380# a_1560_8562# m1_2468_8380# m1_1892_8380# a_182_8562#
+ m1_1508_8380# m1_514_8998# a_1560_9180# m1_322_8140# m1_2180_8140# m1_2372_8998#
+ m1_1988_8140# m1_994_8758# a_182_9180# m1_802_8380# m1_418_8380# m1_1892_8758# VSUBS
+ m1_2276_8380# m1_2468_8758# m1_1700_8380# m1_1508_8758# m1_322_8998# m1_898_8140#
+ m1_130_8140# m1_2180_8998# m1_1796_8140# m1_1090_8140# m1_1988_8998#
Xsky130_fd_pr__nfet_01v8_lvt_324MKY_0 m1_322_8140# m1_610_8758# a_182_9180# m1_994_8380#
+ a_182_8562# a_182_8562# m1_1090_8998# a_182_8562# a_182_8562# a_182_8562# m1_418_8758#
+ m1_226_8380# a_182_8562# a_182_9180# m1_706_8998# a_182_9180# m1_706_8140# m1_514_8140#
+ m1_802_8380# a_182_8562# m1_898_8998# a_182_8562# m1_226_8758# m1_418_8380# a_182_9180#
+ a_182_9180# a_182_9180# a_182_9180# m1_514_8998# a_182_8562# m1_130_8140# m1_1186_8758#
+ m1_1090_8140# m1_610_8380# m1_802_8758# m1_130_8998# m1_322_8998# a_182_9180# m1_1186_8380#
+ a_182_9180# a_182_8562# VSUBS a_182_8562# a_182_9180# m1_994_8758# a_182_9180# m1_898_8140#
+ sky130_fd_pr__nfet_01v8_lvt_324MKY
Xsky130_fd_pr__nfet_01v8_lvt_324MKY_2 m1_2372_8140# m1_2084_8758# a_1560_9180# m1_1700_8380#
+ a_1560_8562# a_1560_8562# m1_1604_8998# a_1560_8562# a_1560_8562# a_1560_8562# m1_2276_8758#
+ m1_2468_8380# a_1560_8562# a_1560_9180# m1_1988_8998# a_1560_9180# m1_1988_8140#
+ m1_2180_8140# m1_1892_8380# a_1560_8562# m1_1796_8998# a_1560_8562# m1_2468_8758#
+ m1_2276_8380# a_1560_9180# a_1560_9180# a_1560_9180# a_1560_9180# m1_2180_8998#
+ a_1560_8562# m1_2564_8140# m1_1508_8758# m1_1604_8140# m1_2084_8380# m1_1892_8758#
+ m1_2564_8998# m1_2372_8998# a_1560_9180# m1_1508_8380# a_1560_9180# a_1560_8562#
+ VSUBS a_1560_8562# a_1560_9180# m1_1700_8758# a_1560_9180# m1_1796_8140# sky130_fd_pr__nfet_01v8_lvt_324MKY
.ends

.subckt sky130_fd_pr__nfet_01v8_ED72KE a_n129_109# a_n753_n1215# a_n753_21# a_n129_727#
+ a_n369_21# a_n705_n509# a_n177_n1215# a_n465_n597# a_255_n509# a_n561_n1215# a_495_n705#
+ a_n609_727# a_n609_109# a_15_1149# a_n273_639# a_399_21# a_n561_1149# a_n81_531#
+ a_447_109# a_447_727# a_399_n1215# a_n177_1149# a_351_n509# a_n417_n509# a_n657_n705#
+ a_n177_n87# a_591_n1215# a_n321_109# a_111_n597# a_n321_727# a_63_n1127# a_n273_531#
+ a_n273_n597# a_n513_n509# a_n797_n1127# a_n33_n1127# a_n129_n509# a_n899_n1301#
+ a_n609_n1127# a_159_109# a_303_n705# a_159_727# a_63_n509# a_n705_n1127# a_n417_n1127#
+ a_n129_n1127# a_n465_639# a_n513_n1127# a_n225_n1127# a_639_727# a_639_109# a_n321_n1127#
+ a_n369_n87# a_n225_n509# a_n465_n705# a_n513_109# a_n513_727# a_687_n597# a_639_n1127#
+ a_n465_531# a_159_n1127# a_447_n1127# a_735_n1127# a_255_n1127# a_543_n1127# a_351_n1127#
+ a_351_727# a_351_109# a_n797_n509# a_n321_n509# a_n33_109# a_n33_727# a_399_1149#
+ a_n81_n597# a_n657_639# a_639_n509# a_111_n705# a_n561_n87# a_n797_727# a_n797_109#
+ a_n225_109# a_n225_727# a_495_639# a_n273_n705# a_15_n1215# a_n705_727# a_n561_21#
+ a_n705_109# a_111_639# a_n177_21# a_n33_n509# a_735_n509# a_n657_531# a_495_n597#
+ a_207_21# a_399_n87# a_543_109# a_543_727# a_591_21# a_495_531# a_111_531# a_591_1149#
+ a_63_727# a_63_109# a_n753_n87# a_n657_n597# a_447_n509# a_687_n705# a_15_n87# a_15_21#
+ a_207_1149# a_n417_109# a_n417_727# a_687_639# a_591_n87# a_303_639# a_n753_1149#
+ a_207_n1215# a_n369_1149# a_255_109# a_255_727# a_543_n509# a_n609_n509# a_159_n509#
+ a_n81_n705# a_207_n87# a_735_727# a_735_109# a_303_n597# a_687_531# a_303_531# a_n369_n1215#
+ a_n81_639#
X0 a_n129_n509# a_n177_n87# a_n225_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X1 a_n321_n1127# a_n369_n1215# a_n417_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X2 a_n417_n509# a_n465_n597# a_n513_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3 a_639_n509# a_591_n87# a_543_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X4 a_n705_n509# a_n753_n87# a_n797_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X5 a_n33_727# a_n81_639# a_n129_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X6 a_351_727# a_303_639# a_255_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X7 a_159_727# a_111_639# a_63_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X8 a_255_727# a_207_1149# a_159_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 a_447_727# a_399_1149# a_351_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X10 a_543_727# a_495_639# a_447_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X11 a_735_727# a_687_639# a_639_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X12 a_63_n1127# a_15_n1215# a_n33_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X13 a_159_n1127# a_111_n705# a_63_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X14 a_639_727# a_591_1149# a_543_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 a_639_n1127# a_591_n1215# a_543_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X16 a_n33_109# a_n81_531# a_n129_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17 a_n33_n509# a_n81_n597# a_n129_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X18 a_351_n509# a_303_n597# a_255_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X19 a_n321_727# a_n369_1149# a_n417_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X20 a_255_n1127# a_207_n1215# a_159_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X21 a_n705_727# a_n753_1149# a_n797_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X22 a_n513_727# a_n561_1149# a_n609_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X23 a_n417_727# a_n465_639# a_n513_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 a_n225_727# a_n273_639# a_n321_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X25 a_n129_727# a_n177_1149# a_n225_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 a_255_109# a_207_21# a_159_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X27 a_351_109# a_303_531# a_255_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X28 a_543_109# a_495_531# a_447_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X29 a_n609_n509# a_n657_n597# a_n705_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X30 a_n417_n1127# a_n465_n705# a_n513_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X31 a_735_n1127# a_687_n705# a_639_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X32 a_n609_727# a_n657_639# a_n705_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 a_159_109# a_111_531# a_63_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X34 a_447_109# a_399_21# a_351_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 a_639_109# a_591_21# a_543_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X36 a_735_109# a_687_531# a_639_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X37 a_n513_n1127# a_n561_n1215# a_n609_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X38 a_351_n1127# a_303_n705# a_255_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X39 a_n513_109# a_n561_21# a_n609_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X40 a_n321_109# a_n369_21# a_n417_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X41 a_n225_109# a_n273_531# a_n321_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X42 a_n705_109# a_n753_21# a_n797_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X43 a_n609_109# a_n657_531# a_n705_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 a_n417_109# a_n465_531# a_n513_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X45 a_n129_109# a_n177_21# a_n225_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 a_255_n509# a_207_n87# a_159_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X47 a_n321_n509# a_n369_n87# a_n417_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X48 a_63_727# a_15_1149# a_n33_727# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X49 a_543_n509# a_495_n597# a_447_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X50 a_n33_n1127# a_n81_n705# a_n129_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X51 a_63_109# a_15_21# a_n33_109# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 a_159_n509# a_111_n597# a_63_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X53 a_n225_n509# a_n273_n597# a_n321_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 a_447_n509# a_399_n87# a_351_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 a_n129_n1127# a_n177_n1215# a_n225_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X56 a_447_n1127# a_399_n1215# a_351_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X57 a_n609_n1127# a_n657_n705# a_n705_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X58 a_n513_n509# a_n561_n87# a_n609_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X59 a_63_n509# a_15_n87# a_n33_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X60 a_735_n509# a_687_n597# a_639_n509# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
X61 a_n225_n1127# a_n273_n705# a_n321_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 a_543_n1127# a_495_n705# a_447_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 a_n705_n1127# a_n753_n1215# a_n797_n1127# a_n899_n1301# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_A574RZ a_761_1345# a_1235_109# a_1235_727# a_n1135_727#
+ a_n1135_109# a_n1135_n1127# a_n1135_n1745# a_n977_n2363# a_n29_n509# a_n503_n1127#
+ a_n503_n1745# a_n129_n2451# a_n29_1963# a_29_n597# a_n29_1345# a_977_21# a_n1235_n2451#
+ a_n129_n597# a_187_21# a_n603_n2451# a_n187_n509# a_n345_n1745# a_n603_639# a_n345_n1127#
+ a_187_n597# a_1077_109# a_n977_109# a_1077_727# a_n977_727# a_1135_639# a_n819_n1745#
+ a_n187_1963# a_n819_n1127# a_n187_1345# a_29_n1215# a_29_n1833# a_n1077_n2451# a_503_n2451#
+ a_n445_n2451# a_129_109# a_129_727# a_n187_n1745# a_n445_21# a_29_1257# a_29_1875#
+ a_n187_n1127# a_n919_n2451# a_1135_n2451# a_n1293_n1745# a_n287_n597# a_n129_1875#
+ a_n1293_n1127# a_n819_n509# a_n129_1257# a_n445_639# a_n661_n1745# a_345_n2451#
+ a_819_n597# a_n819_1963# a_n661_n1127# a_n287_n2451# a_977_639# a_n819_1345# a_187_1257#
+ a_187_1875# a_819_n2451# a_n345_n509# a_n1077_n597# a_345_n597# a_n1077_21# a_n345_1345#
+ a_n345_1963# a_n29_727# a_n761_n2451# a_n29_109# a_187_n2451# a_n1135_n509# a_n919_n597#
+ a_345_21# a_29_21# a_n977_n1127# a_n977_n1745# a_n287_1875# a_n977_n509# a_n287_1257#
+ a_n287_639# a_n1135_1345# a_n1135_1963# a_977_n597# a_n503_727# a_n129_n1215# a_n129_n1833#
+ a_129_n2363# a_n445_n597# a_n503_109# a_819_1257# a_n977_1963# a_819_1875# a_661_n2451#
+ a_603_109# a_603_727# a_n977_1345# a_n1235_n1833# a_n1077_1257# a_n1077_1875# a_n1235_n1215#
+ a_29_639# a_345_1875# a_345_1257# a_n603_n1215# a_n603_n1833# a_603_n2363# a_n1235_n597#
+ a_n603_21# a_n503_n509# a_129_n509# a_n1293_n509# a_n1293_109# a_n1293_727# a_1235_n2363#
+ a_503_n597# a_n919_1875# a_977_n2451# a_n503_1345# a_n919_1257# a_n503_1963# a_n1077_n1833#
+ a_n1077_n1215# a_129_1345# a_129_1963# a_n1293_1963# a_n1293_1345# a_n345_727# a_n919_639#
+ a_503_n1215# a_n445_n1833# a_503_n1833# a_445_n2363# a_n345_109# a_977_1257# a_977_1875#
+ a_n445_n1215# a_445_109# a_445_727# a_503_639# a_n445_1257# a_n445_1875# a_n919_n1833#
+ a_919_n2363# a_n919_n1215# a_n1235_21# a_1135_n1215# a_1135_n1833# a_1077_n2363#
+ a_n603_n597# a_1135_n597# a_n661_n509# a_n761_639# a_287_n509# a_n1235_1257# a_n1235_1875#
+ a_345_n1215# a_n287_n1833# a_345_n1833# a_287_n2363# a_661_n597# a_503_21# a_n287_n1215#
+ a_819_n1833# a_n661_1963# a_503_1875# a_819_n1215# a_n661_1345# a_503_1257# a_287_1963#
+ a_287_1345# a_n187_109# a_n187_727# a_287_727# a_n761_n1833# a_761_n2363# a_287_109#
+ a_345_639# a_n761_n1215# a_187_n1833# a_n29_n2363# a_187_n1215# a_n761_n597# a_n603_1257#
+ a_1135_1875# a_n603_1875# a_919_n509# a_1135_1257# a_129_n1745# a_1135_21# a_n1395_n2537#
+ a_129_n1127# a_661_n1833# a_661_n1215# a_n919_21# a_661_1257# a_919_1963# a_661_1875#
+ a_919_1345# a_n761_21# a_445_n509# a_n129_21# a_n819_727# a_603_n1745# a_n819_109#
+ a_187_639# a_603_n1127# a_n1135_n2363# a_919_109# a_919_727# a_445_1963# a_445_1345#
+ a_1235_n1745# a_977_n1215# a_1235_n1127# a_977_n1833# a_n503_n2363# a_n761_1875#
+ a_n761_1257# a_n1235_639# a_n661_109# a_n661_727# a_445_n1745# a_1077_n509# a_761_727#
+ a_445_n1127# a_761_109# a_919_n1127# a_919_n1745# a_819_21# a_1077_1963# a_1077_n1127#
+ a_1077_n1745# a_661_21# a_1077_1345# a_n345_n2363# a_n819_n2363# a_819_639# a_29_n2451#
+ a_287_n1127# a_287_n1745# a_603_n509# a_603_1345# a_603_1963# a_n187_n2363# a_n1077_639#
+ a_661_639# a_761_n1127# a_n29_n1745# a_761_n1745# a_n29_n1127# a_n1293_n2363# a_n129_639#
+ a_n661_n2363# a_1235_n509# a_761_n509# a_1235_1345# a_1235_1963# a_n287_21# a_761_1963#
X0 a_1235_n1745# a_1135_n1833# a_1077_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_n1135_109# a_n1235_21# a_n1293_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2 a_761_n2363# a_661_n2451# a_603_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3 a_n345_n1127# a_n445_n1215# a_n503_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X4 a_n29_1963# a_n129_1875# a_n187_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X5 a_603_1963# a_503_1875# a_445_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X6 a_1235_n509# a_1135_n597# a_1077_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X7 a_n819_727# a_n919_639# a_n977_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X8 a_n1135_n509# a_n1235_n597# a_n1293_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X9 a_n977_1345# a_n1077_1257# a_n1135_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X10 a_603_n1745# a_503_n1833# a_445_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X11 a_n345_727# a_n445_639# a_n503_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X12 a_1077_1345# a_977_1257# a_919_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X13 a_n661_109# a_n761_21# a_n819_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X14 a_n503_1345# a_n603_1257# a_n661_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X15 a_n819_n1127# a_n919_n1215# a_n977_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X16 a_129_109# a_29_21# a_n29_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X17 a_761_n1745# a_661_n1833# a_603_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X18 a_n977_n1127# a_n1077_n1215# a_n1135_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X19 a_1235_1963# a_1135_1875# a_1077_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X20 a_n503_727# a_n603_639# a_n661_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X21 a_n1135_1963# a_n1235_1875# a_n1293_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X22 a_1235_n1127# a_1135_n1215# a_1077_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X23 a_n187_109# a_n287_21# a_n345_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X24 a_n503_n2363# a_n603_n2451# a_n661_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X25 a_n29_1345# a_n129_1257# a_n187_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X26 a_603_1345# a_503_1257# a_445_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X27 a_287_n2363# a_187_n2451# a_129_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X28 a_n29_727# a_n129_639# a_n187_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X29 a_n819_109# a_n919_21# a_n977_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X30 a_603_n1127# a_503_n1215# a_445_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X31 a_n345_109# a_n445_21# a_n503_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X32 a_n661_n2363# a_n761_n2451# a_n819_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X33 a_n503_n1745# a_n603_n1833# a_n661_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X34 a_761_n1127# a_661_n1215# a_603_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X35 a_n1135_n2363# a_n1235_n2451# a_n1293_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X36 a_n503_109# a_n603_21# a_n661_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X37 a_1077_727# a_977_639# a_919_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X38 a_n1135_1345# a_n1235_1257# a_n1293_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X39 a_1235_1345# a_1135_1257# a_1077_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X40 a_287_n1745# a_187_n1833# a_129_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X41 a_n819_n509# a_n919_n597# a_n977_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X42 a_n661_n1745# a_n761_n1833# a_n819_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X43 a_n29_109# a_n129_21# a_n187_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X44 a_n661_n509# a_n761_n597# a_n819_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X45 a_n29_n2363# a_n129_n2451# a_n187_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X46 a_761_727# a_661_639# a_603_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X47 a_n1135_n1745# a_n1235_n1833# a_n1293_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X48 a_n819_1963# a_n919_1875# a_n977_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X49 a_919_n509# a_819_n597# a_761_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X50 a_n187_n2363# a_n287_n2451# a_n345_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X51 a_n503_n1127# a_n603_n1215# a_n661_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X52 a_287_727# a_187_639# a_129_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X53 a_761_n509# a_661_n597# a_603_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X54 a_1077_109# a_977_21# a_919_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X55 a_n661_1963# a_n761_1875# a_n819_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X56 a_n187_n509# a_n287_n597# a_n345_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X57 a_1235_727# a_1135_639# a_1077_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X58 a_287_n1127# a_187_n1215# a_129_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X59 a_n29_n1745# a_n129_n1833# a_n187_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X60 a_n661_n1127# a_n761_n1215# a_n819_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X61 a_919_727# a_819_639# a_761_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X62 a_919_1963# a_819_1875# a_761_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X63 a_445_727# a_345_639# a_287_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X64 a_n187_n1745# a_n287_n1833# a_n345_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X65 a_n187_1963# a_n287_1875# a_n345_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X66 a_761_1963# a_661_1875# a_603_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X67 a_287_n509# a_187_n597# a_129_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X68 a_761_109# a_661_21# a_603_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X69 a_129_n2363# a_29_n2451# a_n29_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X70 a_n1135_n1127# a_n1235_n1215# a_n1293_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X71 a_n819_1345# a_n919_1257# a_n977_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X72 a_603_727# a_503_639# a_445_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X73 a_287_109# a_187_21# a_129_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X74 a_n661_1345# a_n761_1257# a_n819_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X75 a_1235_109# a_1135_21# a_1077_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X76 a_445_n2363# a_345_n2451# a_287_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X77 a_n29_n1127# a_n129_n1215# a_n187_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X78 a_287_1963# a_187_1875# a_129_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X79 a_129_n1745# a_29_n1833# a_n29_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X80 a_919_1345# a_819_1257# a_761_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X81 a_919_109# a_819_21# a_761_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X82 a_445_109# a_345_21# a_287_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X83 a_n187_n1127# a_n287_n1215# a_n345_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X84 a_n345_n509# a_n445_n597# a_n503_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X85 a_n187_1345# a_n287_1257# a_n345_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X86 a_761_1345# a_661_1257# a_603_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X87 a_919_n2363# a_819_n2451# a_761_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X88 a_445_n1745# a_345_n1833# a_287_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X89 a_129_n509# a_29_n597# a_n29_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X90 a_603_109# a_503_21# a_445_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X91 a_1077_n2363# a_977_n2451# a_919_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X92 a_445_n509# a_345_n597# a_287_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X93 a_n345_1963# a_n445_1875# a_n503_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X94 a_287_1345# a_187_1257# a_129_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X95 a_129_n1127# a_29_n1215# a_n29_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X96 a_919_n1745# a_819_n1833# a_761_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X97 a_129_1963# a_29_1875# a_n29_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X98 a_n345_n2363# a_n445_n2451# a_n503_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X99 a_n977_727# a_n1077_639# a_n1135_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X100 a_1077_n1745# a_977_n1833# a_919_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X101 a_445_1963# a_345_1875# a_287_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X102 a_445_n1127# a_345_n1215# a_287_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X103 a_n977_n509# a_n1077_n597# a_n1135_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X104 a_1077_n509# a_977_n597# a_919_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X105 a_n1135_727# a_n1235_639# a_n1293_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X106 a_n819_n2363# a_n919_n2451# a_n977_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X107 a_n345_1345# a_n445_1257# a_n503_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X108 a_n503_n509# a_n603_n597# a_n661_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X109 a_n345_n1745# a_n445_n1833# a_n503_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X110 a_n977_n2363# a_n1077_n2451# a_n1135_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X111 a_919_n1127# a_819_n1215# a_761_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X112 a_1235_n2363# a_1135_n2451# a_1077_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X113 a_n977_1963# a_n1077_1875# a_n1135_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X114 a_129_1345# a_29_1257# a_n29_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X115 a_n977_109# a_n1077_21# a_n1135_109# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X116 a_1077_1963# a_977_1875# a_919_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X117 a_n661_727# a_n761_639# a_n819_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X118 a_n503_1963# a_n603_1875# a_n661_1963# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X119 a_1077_n1127# a_977_n1215# a_919_n1127# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X120 a_603_n509# a_503_n597# a_445_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X121 a_n29_n509# a_n129_n597# a_n187_n509# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X122 a_445_1345# a_345_1257# a_287_1345# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X123 a_n819_n1745# a_n919_n1833# a_n977_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X124 a_129_727# a_29_639# a_n29_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X125 a_603_n2363# a_503_n2451# a_445_n2363# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X126 a_n977_n1745# a_n1077_n1833# a_n1135_n1745# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X127 a_n187_727# a_n287_639# a_n345_727# a_n1395_n2537# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
.ends

.subckt outd_cmirror_transistors sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n1745# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n2363#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_1345#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n2363#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_21#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n597#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_1257# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n1745#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_1875#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n2363# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_1345# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n2451#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n2451#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n2451#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_1963#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_1345# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n1833# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_1875#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_1875# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_1875# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n1127#
+ a_2_2306# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n2363#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_1963#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n1215# a_2_1688# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_109# a_2_n58# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_1875#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_1345#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_1257# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n1833#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n597# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n1745# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_639#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n2363#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_n509#
+ VSUBS a_2_560# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n1833#
Xsky130_fd_pr__nfet_01v8_ED72KE_0 sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_109# a_2_n58#
+ a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_727# a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_n509#
+ a_2_n58# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_n509# a_2_n58# a_2_n58#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_109#
+ a_2_2306# a_2_2306# a_2_1688# a_2_2306# a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_727# a_2_n58# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_n509# a_2_n58# a_2_560# a_2_n58# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_109#
+ a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_n1127#
+ a_2_1688# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_n509#
+ VSUBS sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_109#
+ a_2_n58# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n129_n1127# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_n1127#
+ a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_n509# a_2_n58# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n513_727# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_n1127#
+ a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_n1127# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_n1127#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_351_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n321_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_727#
+ a_2_2306# a_2_560# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_639_n509# a_2_n58#
+ a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_727# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n797_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n225_727#
+ a_2_2306# a_2_n58# a_2_n58# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_727# a_2_1688#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n705_109# a_2_2306# a_2_1688# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n33_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_n509# a_2_1688# a_2_560# a_2_1688# a_2_560#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_727#
+ a_2_1688# a_2_1688# a_2_1688# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_63_109# a_2_560# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_447_n509#
+ a_2_n58# a_2_560# a_2_1688# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_109#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_n417_727# a_2_2306# a_2_560# a_2_2306# a_2_2306#
+ a_2_n58# a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_109# sky130_fd_pr__nfet_01v8_ED72KE_0/a_255_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_543_n509# sky130_fd_pr__nfet_01v8_ED72KE_0/a_n609_n509#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_159_n509# a_2_n58# a_2_560# sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_727#
+ sky130_fd_pr__nfet_01v8_ED72KE_0/a_735_109# a_2_560# a_2_1688# a_2_1688# a_2_n58#
+ a_2_2306# sky130_fd_pr__nfet_01v8_ED72KE
Xsky130_fd_pr__nfet_01v8_A574RZ_0 sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n2451#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n977_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n445_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_n597# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_503_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_109#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_345_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_n1215# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_n597#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n603_1875# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1135_21# VSUBS sky130_fd_pr__nfet_01v8_A574RZ_0/a_129_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n1833# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n919_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_1257#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_187_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1135_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_1345#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n1215#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_977_n1833#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n503_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_1875#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n761_1257# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1235_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_727#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_727# sky130_fd_pr__nfet_01v8_A574RZ_0/a_445_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_109# sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_919_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_1963# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_21#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1077_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n345_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n819_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_819_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_29_n2451# sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_287_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_603_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n187_n2363# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1077_639#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_661_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n1127#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n1745# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n1745#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n29_n1127# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n1293_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n129_639# sky130_fd_pr__nfet_01v8_A574RZ_0/a_n661_n2363#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_n509# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_n509#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_1345# sky130_fd_pr__nfet_01v8_A574RZ_0/a_1235_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ_0/a_n287_21# sky130_fd_pr__nfet_01v8_A574RZ_0/a_761_1963#
+ sky130_fd_pr__nfet_01v8_A574RZ
.ends

.subckt outd_cmirror_64t m1_220_5610# m1_0_80# m1_130_5370# VSUBS
Xoutd_cmirror_transistors_0 m1_220_5610# m1_130_5370# m1_130_5370# m1_220_5610# m1_130_5370#
+ VSUBS m1_130_5370# VSUBS m1_220_5610# VSUBS m1_0_80# m1_0_80# VSUBS VSUBS VSUBS
+ m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_220_5610# m1_130_5370# m1_220_5610# m1_220_5610#
+ m1_220_5610# m1_0_80# m1_220_5610# m1_130_5370# m1_220_5610# m1_220_5610# m1_220_5610#
+ VSUBS VSUBS m1_220_5610# VSUBS m1_220_5610# m1_0_80# VSUBS VSUBS m1_0_80# m1_0_80#
+ m1_220_5610# m1_0_80# m1_130_5370# m1_220_5610# m1_220_5610# m1_220_5610# m1_0_80#
+ m1_220_5610# m1_0_80# m1_220_5610# m1_220_5610# m1_220_5610# m1_0_80# m1_220_5610#
+ m1_0_80# m1_220_5610# m1_220_5610# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# VSUBS
+ VSUBS VSUBS m1_130_5370# m1_220_5610# m1_130_5370# VSUBS VSUBS m1_220_5610# m1_0_80#
+ VSUBS VSUBS m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_130_5370# m1_0_80# VSUBS
+ VSUBS m1_220_5610# m1_130_5370# VSUBS m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610#
+ m1_0_80# m1_0_80# VSUBS VSUBS m1_0_80# VSUBS VSUBS m1_220_5610# m1_220_5610# m1_220_5610#
+ m1_130_5370# m1_220_5610# m1_130_5370# m1_130_5370# m1_220_5610# m1_220_5610# m1_0_80#
+ m1_130_5370# m1_220_5610# m1_220_5610# VSUBS VSUBS VSUBS m1_220_5610# m1_220_5610#
+ m1_220_5610# m1_130_5370# m1_220_5610# m1_0_80# m1_130_5370# m1_220_5610# m1_0_80#
+ m1_0_80# VSUBS m1_130_5370# VSUBS VSUBS m1_130_5370# m1_220_5610# m1_220_5610# m1_0_80#
+ m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_220_5610# m1_220_5610# m1_0_80# VSUBS
+ m1_220_5610# m1_0_80# VSUBS m1_0_80# m1_0_80# VSUBS VSUBS m1_220_5610# m1_0_80#
+ m1_0_80# m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS VSUBS m1_0_80# m1_0_80# m1_220_5610#
+ m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS m1_220_5610#
+ VSUBS m1_220_5610# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS
+ m1_220_5610# m1_130_5370# m1_130_5370# m1_0_80# VSUBS VSUBS VSUBS VSUBS m1_220_5610#
+ m1_0_80# m1_220_5610# m1_130_5370# m1_0_80# m1_130_5370# m1_0_80# m1_220_5610# m1_0_80#
+ VSUBS m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_220_5610# m1_220_5610# m1_0_80# m1_0_80#
+ m1_0_80# m1_0_80# m1_0_80# m1_130_5370# m1_130_5370# m1_130_5370# m1_0_80# m1_0_80#
+ m1_0_80# m1_0_80# m1_0_80# m1_130_5370# m1_0_80# m1_0_80# m1_220_5610# m1_220_5610#
+ m1_220_5610# VSUBS m1_220_5610# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_0_80#
+ VSUBS m1_220_5610# m1_0_80# m1_0_80# VSUBS m1_220_5610# VSUBS m1_0_80# m1_0_80#
+ VSUBS VSUBS m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80#
+ m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_220_5610#
+ m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# m1_0_80#
+ m1_220_5610# m1_220_5610# m1_220_5610# m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS m1_220_5610#
+ m1_130_5370# m1_130_5370# m1_220_5610# m1_0_80# m1_0_80# m1_130_5370# m1_130_5370#
+ m1_220_5610# m1_0_80# m1_0_80# m1_130_5370# m1_0_80# m1_0_80# m1_130_5370# VSUBS
+ m1_220_5610# m1_220_5610# VSUBS VSUBS m1_130_5370# m1_0_80# VSUBS m1_0_80# VSUBS
+ m1_0_80# VSUBS m1_130_5370# m1_0_80# m1_130_5370# m1_220_5610# m1_0_80# m1_220_5610#
+ VSUBS VSUBS m1_0_80# VSUBS VSUBS m1_220_5610# m1_0_80# m1_220_5610# m1_0_80# m1_0_80#
+ VSUBS m1_0_80# m1_0_80# m1_0_80# VSUBS VSUBS VSUBS VSUBS VSUBS m1_220_5610# m1_220_5610#
+ m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610# m1_220_5610#
+ VSUBS m1_0_80# m1_0_80# m1_0_80# m1_0_80# m1_0_80# outd_cmirror_transistors
.ends

.subckt outd_stage2 m1_370_11400# m1_2350_11400# outd_cmirror_64t_4/m1_0_80# dw_60_8030#
+ m1_1850_8370# m2_7240_7300# cmirror_out m1_250_8900# VN
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_0 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_1 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_2 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_3 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_4 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_5 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_6 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_8 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_7 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_9 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_10 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_11 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_12 m1_2350_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_13 m1_370_11400# dw_60_8030# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_14 dw_60_8030# m1_370_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xsky130_fd_pr__res_high_po_5p73_PA2QZX_15 dw_60_8030# m1_2350_11400# VN sky130_fd_pr__res_high_po_5p73_PA2QZX
Xoutd_diffamp_0 cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_370_11400# m1_2350_11400# m1_2350_11400# cmirror_out cmirror_out cmirror_out
+ cmirror_out m1_370_11400# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400#
+ cmirror_out m1_1850_8370# cmirror_out cmirror_out m1_250_8900# cmirror_out m1_370_11400#
+ m1_1850_8370# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400# cmirror_out
+ m1_250_8900# cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_2350_11400# m1_370_11400# m1_2350_11400# outd_diffamp
Xoutd_cmirror_64t_0 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
Xoutd_diffamp_1 cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_370_11400# m1_2350_11400# m1_2350_11400# cmirror_out cmirror_out cmirror_out
+ cmirror_out m1_370_11400# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400#
+ cmirror_out m1_1850_8370# cmirror_out cmirror_out m1_250_8900# cmirror_out m1_370_11400#
+ m1_1850_8370# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400# cmirror_out
+ m1_250_8900# cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_2350_11400# m1_370_11400# m1_2350_11400# outd_diffamp
Xoutd_cmirror_64t_2 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
Xoutd_cmirror_64t_1 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
Xoutd_diffamp_2 cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_370_11400# m1_2350_11400# m1_2350_11400# cmirror_out cmirror_out cmirror_out
+ cmirror_out m1_370_11400# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400#
+ cmirror_out m1_1850_8370# cmirror_out cmirror_out m1_250_8900# cmirror_out m1_370_11400#
+ m1_1850_8370# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400# cmirror_out
+ m1_250_8900# cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_2350_11400# m1_370_11400# m1_2350_11400# outd_diffamp
Xoutd_cmirror_64t_3 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
Xoutd_diffamp_3 cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_370_11400# m1_2350_11400# m1_2350_11400# cmirror_out cmirror_out cmirror_out
+ cmirror_out m1_370_11400# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400#
+ cmirror_out m1_1850_8370# cmirror_out cmirror_out m1_250_8900# cmirror_out m1_370_11400#
+ m1_1850_8370# m1_370_11400# m1_2350_11400# m1_2350_11400# m1_2350_11400# cmirror_out
+ m1_250_8900# cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out cmirror_out
+ cmirror_out cmirror_out m1_370_11400# m1_370_11400# m1_370_11400# m1_2350_11400#
+ m1_2350_11400# m1_370_11400# m1_2350_11400# outd_diffamp
Xoutd_cmirror_64t_4 m2_7240_7300# outd_cmirror_64t_4/m1_0_80# cmirror_out VN outd_cmirror_64t
.ends

.subckt sky130_fd_pr__nfet_01v8_DJG2KN a_n29_n509# a_29_n597# a_n187_n509# a_n129_n597#
+ a_129_109# a_n289_n683# a_n29_109# a_29_21# a_129_n509# a_n187_109# a_n129_21#
X0 a_129_109# a_29_21# a_n29_109# a_n289_n683# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_n29_109# a_n129_21# a_n187_109# a_n289_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2 a_129_n509# a_29_n597# a_n29_n509# a_n289_n683# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3 a_n29_n509# a_n129_n597# a_n187_n509# a_n289_n683# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt outd_stage3 m4_40470_12200# m3_11690_14240# m2_40400_9110# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ outd_stage2_3/cmirror_out m4_40470_12880# m2_40400_10380# VSUBS
Xoutd_stage2_0 m4_40470_12880# m4_40470_12200# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ m3_11690_14240# m2_40400_9110# m2_41490_8160# outd_stage2_3/cmirror_out m2_40400_10380#
+ VSUBS outd_stage2
Xoutd_stage2_1 m4_40470_12880# m4_40470_12200# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ m3_11690_14240# m2_40400_9110# m2_41490_8160# outd_stage2_3/cmirror_out m2_40400_10380#
+ VSUBS outd_stage2
Xoutd_stage2_2 m4_40470_12880# m4_40470_12200# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ m3_11690_14240# m2_40400_9110# m2_41490_8160# outd_stage2_3/cmirror_out m2_40400_10380#
+ VSUBS outd_stage2
Xoutd_stage2_3 m4_40470_12880# m4_40470_12200# outd_stage2_3/outd_cmirror_64t_4/m1_0_80#
+ m3_11690_14240# m2_40400_9110# m2_41490_8160# outd_stage2_3/cmirror_out m2_40400_10380#
+ VSUBS outd_stage2
.ends

.subckt sky130_fd_pr__nfet_01v8_LH2JGW a_n81_n288# a_63_n200# a_n33_n200# a_15_222#
+ a_n227_n374# a_n125_n200#
X0 a_n33_n200# a_n81_n288# a_n125_n200# a_n227_n374# sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X1 a_63_n200# a_15_222# a_n33_n200# a_n227_n374# sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__res_high_po_2p85_8GE2XM a_n1512_n1032# a_n694_n1032# a_124_n1032#
+ a_n1512_600# a_n1642_n1162# a_942_n1032# a_124_600# a_942_600# a_n694_600#
X0 a_n1512_n1032# a_n1512_600# a_n1642_n1162# sky130_fd_pr__res_high_po_2p85 l=6e+06u
X1 a_n694_n1032# a_n694_600# a_n1642_n1162# sky130_fd_pr__res_high_po_2p85 l=6e+06u
X2 a_942_n1032# a_942_600# a_n1642_n1162# sky130_fd_pr__res_high_po_2p85 l=6e+06u
X3 a_124_n1032# a_124_600# a_n1642_n1162# sky130_fd_pr__res_high_po_2p85 l=6e+06u
.ends

.subckt outd_stage1 outd_cmirror_64t_0/m1_0_80# m1_n1500_10180# m1_1860_8350# isource_out
+ m1_1830_10170# m1_260_8900# dw_70_8020# VN
Xoutd_cmirror_64t_0 outd_cmirror_64t_0/m1_220_5610# outd_cmirror_64t_0/m1_0_80# isource_out
+ VN outd_cmirror_64t
Xoutd_diffamp_0 isource_out isource_out isource_out isource_out isource_out isource_out
+ isource_out isource_out m1_n1500_10180# m1_n1500_10180# m1_n1500_10180# m1_1830_10170#
+ m1_n1500_10180# m1_1830_10170# m1_1830_10170# isource_out isource_out isource_out
+ isource_out m1_n1500_10180# m1_n1500_10180# m1_1830_10170# m1_1830_10170# m1_1830_10170#
+ isource_out m1_1860_8350# isource_out isource_out m1_260_8900# isource_out m1_n1500_10180#
+ m1_1860_8350# m1_n1500_10180# m1_1830_10170# m1_1830_10170# m1_1830_10170# isource_out
+ m1_260_8900# isource_out isource_out isource_out isource_out isource_out isource_out
+ isource_out isource_out m1_n1500_10180# m1_n1500_10180# m1_n1500_10180# m1_1830_10170#
+ m1_1830_10170# m1_n1500_10180# m1_1830_10170# outd_diffamp
Xsky130_fd_pr__res_high_po_2p85_8GE2XM_0 m1_n1500_10180# m1_n1500_10180# m1_n1500_10180#
+ dw_70_8020# VN m1_n1500_10180# dw_70_8020# dw_70_8020# dw_70_8020# sky130_fd_pr__res_high_po_2p85_8GE2XM
Xsky130_fd_pr__res_high_po_2p85_8GE2XM_1 m1_1830_10170# m1_1830_10170# m1_1830_10170#
+ dw_70_8020# VN m1_1830_10170# dw_70_8020# dw_70_8020# dw_70_8020# sky130_fd_pr__res_high_po_2p85_8GE2XM
.ends

.subckt outd
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_6 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_7 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_1_WXTTNJ_0 VN I_Bias sky130_fd_pr__cap_mim_m3_1_WXTTNJ
Xsky130_fd_pr__cap_mim_m3_1_WXTTNJ_1 VN I_Bias sky130_fd_pr__cap_mim_m3_1_WXTTNJ
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_8 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xoutd_stage2_0 V_da2_N V_da2_P I_Bias VP V_da1_P outd_stage2_0/m2_7240_7300# VM1_D
+ V_da1_N VN outd_stage2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_9 VN InputRef sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__nfet_01v8_DJG2KN_0 m1_n19890_7120# I_Bias VN I_Bias VN VN m1_n19890_7120#
+ I_Bias VN VN I_Bias sky130_fd_pr__nfet_01v8_DJG2KN
Xoutd_stage3_0 OutputP VP V_da2_P I_Bias VM14D OutputN V_da2_N VN outd_stage3
Xsky130_fd_pr__nfet_01v8_LH2JGW_0 I_Bias m1_n19890_7120# I_Bias I_Bias VN m1_n19890_7120#
+ sky130_fd_pr__nfet_01v8_LH2JGW
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_10 VN InputRef sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xoutd_stage1_0 I_Bias V_da1_P InputRef outd_stage1_0/isource_out V_da1_N InputSignal
+ VP VN outd_stage1
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_0 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_1 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_2 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_4 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_3 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
Xsky130_fd_pr__cap_mim_m3_2_LJ5JLG_5 VP VN sky130_fd_pr__cap_mim_m3_2_LJ5JLG#2
.ends

