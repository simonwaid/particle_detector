magic
tech sky130A
magscale 1 2
timestamp 1645541123
<< error_p >>
rect -530 291 530 318
rect -530 -318 530 -291
<< nwell >>
rect -633 -291 633 291
<< pwell >>
rect -743 291 743 401
rect -743 -291 -633 291
rect 633 -291 743 291
rect -743 -401 743 -291
<< varactor >>
rect -500 -200 500 200
<< psubdiff >>
rect -707 331 -611 365
rect 611 331 707 365
rect -707 269 -673 331
rect 673 269 707 331
rect -707 -331 -673 -269
rect 673 -331 707 -269
rect -707 -365 -611 -331
rect 611 -365 707 -331
<< nsubdiff >>
rect -597 176 -500 200
rect -597 -176 -585 176
rect -551 -176 -500 176
rect -597 -200 -500 -176
rect 500 176 597 200
rect 500 -176 551 176
rect 585 -176 597 176
rect 500 -200 597 -176
<< psubdiffcont >>
rect -611 331 611 365
rect -707 -269 -673 269
rect 673 -269 707 269
rect -611 -365 611 -331
<< nsubdiffcont >>
rect -585 -176 -551 176
rect 551 -176 585 176
<< poly >>
rect -500 272 500 288
rect -500 238 -484 272
rect 484 238 500 272
rect -500 200 500 238
rect -500 -238 500 -200
rect -500 -272 -484 -238
rect 484 -272 500 -238
rect -500 -288 500 -272
<< polycont >>
rect -484 238 484 272
rect -484 -272 484 -238
<< locali >>
rect -707 331 -611 365
rect 611 331 707 365
rect -707 269 -673 331
rect -500 238 -484 272
rect 484 238 500 272
rect 673 269 707 331
rect -585 176 -551 192
rect -585 -192 -551 -176
rect 551 176 585 192
rect 551 -192 585 -176
rect -707 -331 -673 -269
rect -500 -272 -484 -238
rect 484 -272 500 -238
rect 673 -331 707 -269
rect -707 -365 -611 -331
rect 611 -365 707 -331
<< viali >>
rect -484 238 484 272
rect -585 -176 -551 176
rect 551 -176 585 176
rect -484 -272 484 -238
<< metal1 >>
rect -496 272 496 278
rect -496 238 -484 272
rect 484 238 496 272
rect -496 232 496 238
rect -591 176 -545 188
rect -591 -176 -585 176
rect -551 -176 -545 176
rect -591 -188 -545 -176
rect 545 176 591 188
rect 545 -176 551 176
rect 585 -176 591 176
rect 545 -188 591 -176
rect -496 -238 496 -232
rect -496 -272 -484 -238
rect 484 -272 496 -238
rect -496 -278 496 -272
<< properties >>
string FIXED_BBOX -690 -348 690 348
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 2 l 5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
