magic
tech sky130B
magscale 1 2
timestamp 1654704381
<< metal1 >>
rect 2240 8950 2290 9310
rect 3040 9250 3400 9310
rect 3330 8960 3380 9250
rect 5510 8960 5560 9320
rect 6340 9250 6640 9310
rect 8520 9220 8820 9280
rect 10690 9220 10990 9280
rect 12900 9220 13200 9280
rect 15070 9220 15370 9280
rect 17260 9220 17560 9280
rect 19420 9220 19710 9280
rect 2240 6670 2290 7030
rect 5510 7020 5560 7050
rect 3080 6960 3440 7020
rect 4140 6960 4500 7020
rect 5240 6960 5600 7020
rect 6370 6960 6650 7020
rect 3330 6660 3380 6960
rect 4420 6650 4470 6960
rect 5510 6690 5560 6960
rect 8520 6940 8800 7000
rect 10700 6940 10980 7000
rect 12900 6940 13180 7000
rect 15060 6940 15340 7000
rect 17260 6940 17540 7000
rect 19420 6940 19710 7000
rect 3330 4730 3380 4740
rect 60 4370 110 4720
rect 2240 4370 2290 4730
rect 3070 4670 3430 4730
rect 4120 4670 4480 4730
rect 5270 4670 5630 4730
rect 6360 4670 6650 4730
rect 3330 4380 3380 4670
rect 4420 4370 4470 4670
rect 5510 4360 5560 4670
rect 8520 4660 8830 4720
rect 10680 4660 10990 4720
rect 12880 4660 13190 4720
rect 15040 4660 15350 4720
rect 17260 4660 17570 4720
rect 19410 4660 19700 4720
rect 840 2340 910 2410
rect 1030 2340 1040 2410
rect 1150 2380 5630 2440
rect 6360 2380 6670 2440
rect 8520 2380 8830 2440
rect 10720 2380 11030 2440
rect 12880 2380 13190 2440
rect 15050 2380 15360 2440
rect 17210 2380 17520 2440
rect 19450 2380 19740 2440
rect 1760 2320 1920 2380
rect 1750 2250 1760 2320
rect 1920 2250 1930 2320
rect 5360 2280 5520 2380
rect 640 2160 650 2240
rect 860 2160 870 2240
rect 5350 2190 5360 2280
rect 5520 2190 5530 2280
rect 640 2080 870 2160
rect 920 2070 1200 2120
rect 1990 2070 2280 2120
rect 3040 2070 3330 2120
<< via1 >>
rect 910 2340 1030 2410
rect 1760 2250 1920 2320
rect 650 2160 860 2240
rect 5360 2190 5520 2280
<< metal2 >>
rect 2330 11250 2620 11260
rect 2330 11070 2620 11080
rect 3440 11250 3730 11260
rect 3440 11070 3730 11080
rect 5590 11250 5880 11260
rect 5590 11070 5880 11080
rect 3280 10400 3360 10410
rect 3360 10250 4140 10400
rect 3280 10240 3360 10250
rect 2990 9970 3560 10120
rect 3280 9770 3360 9780
rect 3360 9620 4140 9770
rect 3280 9610 3360 9620
rect 2330 8960 2620 8970
rect 2330 8780 2620 8790
rect 3110 8460 3230 9350
rect 3430 8960 3720 8970
rect 3430 8780 3720 8790
rect 4490 8960 4780 8970
rect 4490 8780 4780 8790
rect 5590 8960 5880 8970
rect 5590 8780 5880 8790
rect 6380 8570 6500 9490
rect 160 6800 430 6810
rect 160 6490 430 6500
rect 2330 6670 2620 6680
rect 2330 6490 2620 6500
rect 3110 6330 3230 7220
rect 3430 6670 3720 6680
rect 3430 6490 3720 6500
rect 4200 6300 4320 7190
rect 4490 6670 4780 6680
rect 4490 6490 4780 6500
rect 5290 6250 5410 7170
rect 5590 6670 5880 6680
rect 5590 6490 5880 6500
rect 6380 6260 6500 7180
rect 160 4520 430 4530
rect 160 4210 430 4220
rect 2330 4370 2620 4380
rect 2330 4190 2620 4200
rect 3110 3920 3230 4810
rect 3430 4380 3720 4390
rect 3430 4200 3720 4210
rect 4200 3920 4320 4810
rect 4490 4380 4780 4390
rect 4490 4200 4780 4210
rect 5290 3930 5410 4850
rect 5590 4380 5880 4390
rect 5590 4200 5880 4210
rect 6380 3850 6500 4770
rect 4310 2460 4530 2640
rect 770 2410 1120 2420
rect 1030 2350 1120 2410
rect 1030 2340 1450 2350
rect 770 2330 1450 2340
rect 1000 2310 1450 2330
rect 650 2240 860 2250
rect 1000 2230 1250 2310
rect 1380 2230 1450 2310
rect 1760 2320 1920 2330
rect 1760 2240 1920 2250
rect 5360 2280 5520 2290
rect 1000 2210 1450 2230
rect 650 2150 860 2160
rect 1330 1980 1450 2210
rect 5360 2180 5520 2190
rect 3220 480 3670 630
rect 390 330 610 340
rect 390 10 610 20
rect 1480 330 1700 340
rect 1480 10 1700 20
rect 2570 330 2790 340
rect 2570 10 2790 20
rect 3660 330 3880 340
rect 3660 10 3880 20
<< via2 >>
rect 2330 11080 2620 11250
rect 3440 11080 3730 11250
rect 5590 11080 5880 11250
rect 3280 10250 3360 10400
rect 3280 9620 3360 9770
rect 2330 8790 2620 8960
rect 3430 8790 3720 8960
rect 4490 8790 4780 8960
rect 5590 8790 5880 8960
rect 160 6500 430 6800
rect 2330 6500 2620 6670
rect 3430 6500 3720 6670
rect 4490 6500 4780 6670
rect 5590 6500 5880 6670
rect 160 4220 430 4520
rect 2330 4200 2620 4370
rect 3430 4210 3720 4380
rect 4490 4210 4780 4380
rect 5590 4210 5880 4380
rect 770 2340 910 2410
rect 910 2340 1030 2410
rect 650 2160 860 2240
rect 1250 2230 1380 2310
rect 1760 2250 1920 2320
rect 5360 2190 5520 2280
rect 390 20 610 330
rect 1480 20 1700 330
rect 2570 20 2790 330
rect 3660 20 3880 330
<< metal3 >>
rect 2330 11410 2620 11430
rect 3430 11410 3720 11430
rect 4490 11410 4780 11430
rect 5590 11410 5880 11430
rect 150 11390 440 11410
rect 150 11020 180 11390
rect 450 11020 460 11390
rect 2320 11080 2330 11410
rect 2620 11080 2630 11410
rect 2320 11075 2630 11080
rect 3430 11080 3440 11410
rect 3730 11080 3740 11410
rect 4480 11080 4490 11410
rect 4780 11080 4790 11410
rect 5580 11080 5590 11410
rect 5880 11080 5890 11410
rect 3430 11075 3740 11080
rect 150 6800 440 11020
rect 2330 8965 2620 11075
rect 3270 10400 3370 10405
rect 3020 10390 3280 10400
rect 2820 10250 3280 10390
rect 3360 10250 3370 10400
rect 2820 9770 3060 10250
rect 3270 10245 3370 10250
rect 3270 9770 3370 9775
rect 2820 9620 3280 9770
rect 3360 9620 3370 9770
rect 2320 8960 2630 8965
rect 2320 8790 2330 8960
rect 2620 8790 2630 8960
rect 2320 8785 2630 8790
rect 150 6500 160 6800
rect 430 6500 440 6800
rect 2330 6675 2620 8785
rect 150 4520 440 6500
rect 2320 6670 2630 6675
rect 2320 6500 2330 6670
rect 2620 6500 2630 6670
rect 2320 6495 2630 6500
rect 660 5220 790 5350
rect 150 4220 160 4520
rect 430 4220 440 4520
rect 2330 4375 2620 6495
rect 150 4210 440 4220
rect 2320 4370 2630 4375
rect 2320 4200 2330 4370
rect 2620 4200 2630 4370
rect 2320 4195 2630 4200
rect 770 2415 1010 2890
rect 760 2410 1040 2415
rect 760 2340 770 2410
rect 1030 2340 1040 2410
rect 760 2335 1040 2340
rect 1730 2370 1970 2880
rect 2820 2760 3060 9620
rect 3270 9615 3370 9620
rect 3430 8965 3720 11075
rect 4490 8965 4780 11080
rect 5580 11075 5890 11080
rect 5590 8965 5880 11075
rect 6690 11050 6700 11380
rect 6990 11050 7000 11380
rect 7780 11050 7790 11380
rect 8080 11050 8090 11380
rect 8870 11050 8880 11380
rect 9170 11050 9180 11380
rect 9960 11050 9970 11380
rect 10260 11050 10270 11380
rect 11050 11050 11060 11380
rect 11350 11050 11360 11380
rect 12140 11050 12150 11380
rect 12440 11050 12450 11380
rect 13230 11050 13240 11380
rect 13530 11050 13540 11380
rect 14320 11050 14330 11380
rect 14620 11050 14630 11380
rect 15410 11050 15420 11380
rect 15710 11050 15720 11380
rect 16500 11050 16510 11380
rect 16800 11050 16810 11380
rect 17590 11050 17600 11380
rect 17890 11050 17900 11380
rect 18680 11050 18690 11380
rect 18980 11050 18990 11380
rect 19770 11050 19780 11380
rect 20070 11050 20080 11380
rect 20860 11050 20870 11380
rect 21160 11050 21170 11380
rect 3420 8960 3730 8965
rect 3420 8790 3430 8960
rect 3720 8790 3730 8960
rect 3420 8785 3730 8790
rect 4480 8960 4790 8965
rect 4480 8790 4490 8960
rect 4780 8790 4790 8960
rect 4480 8785 4790 8790
rect 5580 8960 5890 8965
rect 5580 8790 5590 8960
rect 5880 8790 5890 8960
rect 5580 8785 5890 8790
rect 3430 6675 3720 8785
rect 3420 6670 3730 6675
rect 3420 6500 3430 6670
rect 3720 6500 3730 6670
rect 3420 6495 3730 6500
rect 3430 4385 3720 6495
rect 3420 4380 3730 4385
rect 3420 4210 3430 4380
rect 3720 4210 3730 4380
rect 3420 4205 3730 4210
rect 3430 4200 3720 4205
rect 3900 2970 4140 8100
rect 4490 6675 4780 8785
rect 4480 6670 4790 6675
rect 4480 6500 4490 6670
rect 4780 6500 4790 6670
rect 4480 6495 4790 6500
rect 4490 4385 4780 6495
rect 4480 4380 4790 4385
rect 4480 4210 4490 4380
rect 4780 4210 4790 4380
rect 4480 4205 4790 4210
rect 4490 4200 4780 4205
rect 5000 2970 5240 8100
rect 5590 6675 5880 8785
rect 5580 6670 5890 6675
rect 5580 6500 5590 6670
rect 5880 6500 5890 6670
rect 5580 6495 5890 6500
rect 5590 4385 5880 6495
rect 5580 4380 5890 4385
rect 5580 4210 5590 4380
rect 5880 4210 5890 4380
rect 5580 4205 5890 4210
rect 5590 4200 5880 4205
rect 3900 2760 5240 2970
rect 6090 2760 6330 10390
rect 7560 2710 7750 2890
rect 9720 2720 9900 2870
rect 11910 2730 12060 2850
rect 14070 2720 14220 2840
rect 16330 2720 16470 2820
rect 18470 2730 18610 2830
rect 20660 2760 20840 2850
rect 1730 2320 3070 2370
rect 1240 2310 1390 2315
rect 30 2240 880 2270
rect 30 2160 650 2240
rect 860 2160 880 2240
rect 1240 2230 1250 2310
rect 1380 2230 1390 2310
rect 1240 2225 1390 2230
rect 1730 2250 1760 2320
rect 1920 2250 3070 2320
rect 1730 2200 3070 2250
rect 30 2130 880 2160
rect 640 1910 880 2130
rect 2820 2060 3070 2200
rect 5340 2180 5350 2320
rect 5540 2180 5550 2320
rect 2810 1890 4150 2060
rect 370 340 380 450
rect 100 40 380 340
rect 760 340 770 450
rect 1460 340 1470 450
rect 760 40 1470 340
rect 1850 340 1860 450
rect 2550 340 2560 450
rect 1850 40 2560 340
rect 2940 340 2950 450
rect 3640 340 3650 450
rect 2940 40 3650 340
rect 4030 40 4040 450
rect 100 20 390 40
rect 610 20 1480 40
rect 1700 20 2570 40
rect 2790 20 3660 40
rect 3880 20 3890 40
rect 380 15 620 20
rect 1470 15 1710 20
rect 2560 15 2800 20
rect 3650 15 3890 20
<< via3 >>
rect 180 11020 450 11390
rect 2330 11250 2620 11410
rect 2330 11080 2620 11250
rect 3440 11250 3730 11410
rect 3440 11080 3730 11250
rect 4490 11080 4780 11410
rect 5590 11250 5880 11410
rect 5590 11080 5880 11250
rect 6700 11050 6990 11380
rect 7790 11050 8080 11380
rect 8880 11050 9170 11380
rect 9970 11050 10260 11380
rect 11060 11050 11350 11380
rect 12150 11050 12440 11380
rect 13240 11050 13530 11380
rect 14330 11050 14620 11380
rect 15420 11050 15710 11380
rect 16510 11050 16800 11380
rect 17600 11050 17890 11380
rect 18690 11050 18980 11380
rect 19780 11050 20070 11380
rect 20870 11050 21160 11380
rect 1250 2230 1380 2310
rect 5350 2280 5540 2320
rect 5350 2190 5360 2280
rect 5360 2190 5520 2280
rect 5520 2190 5540 2280
rect 5350 2180 5540 2190
rect 380 330 760 450
rect 380 40 390 330
rect 390 40 610 330
rect 610 40 760 330
rect 1470 330 1850 450
rect 1470 40 1480 330
rect 1480 40 1700 330
rect 1700 40 1850 330
rect 2560 330 2940 450
rect 2560 40 2570 330
rect 2570 40 2790 330
rect 2790 40 2940 330
rect 3650 330 4030 450
rect 3650 40 3660 330
rect 3660 40 3880 330
rect 3880 40 4030 330
<< metal4 >>
rect 2329 11410 2621 11411
rect 179 11390 451 11391
rect 179 11020 180 11390
rect 450 11020 451 11390
rect 2329 11080 2330 11410
rect 2620 11080 2621 11410
rect 2329 11079 2621 11080
rect 3439 11410 3731 11411
rect 3439 11080 3440 11410
rect 3730 11080 3731 11410
rect 3439 11079 3731 11080
rect 4489 11410 4781 11411
rect 4489 11080 4490 11410
rect 4780 11080 4781 11410
rect 4489 11079 4781 11080
rect 5589 11410 5881 11411
rect 5589 11080 5590 11410
rect 5880 11080 5881 11410
rect 5589 11079 5881 11080
rect 6699 11380 6991 11381
rect 6699 11050 6700 11380
rect 6990 11050 6991 11380
rect 6699 11049 6991 11050
rect 7789 11380 8081 11381
rect 7789 11050 7790 11380
rect 8080 11050 8081 11380
rect 7789 11049 8081 11050
rect 8879 11380 9171 11381
rect 8879 11050 8880 11380
rect 9170 11050 9171 11380
rect 8879 11049 9171 11050
rect 9969 11380 10261 11381
rect 9969 11050 9970 11380
rect 10260 11050 10261 11380
rect 9969 11049 10261 11050
rect 11059 11380 11351 11381
rect 11059 11050 11060 11380
rect 11350 11050 11351 11380
rect 11059 11049 11351 11050
rect 12149 11380 12441 11381
rect 12149 11050 12150 11380
rect 12440 11050 12441 11380
rect 12149 11049 12441 11050
rect 13239 11380 13531 11381
rect 13239 11050 13240 11380
rect 13530 11050 13531 11380
rect 13239 11049 13531 11050
rect 14329 11380 14621 11381
rect 14329 11050 14330 11380
rect 14620 11050 14621 11380
rect 14329 11049 14621 11050
rect 15419 11380 15711 11381
rect 15419 11050 15420 11380
rect 15710 11050 15711 11380
rect 15419 11049 15711 11050
rect 16509 11380 16801 11381
rect 16509 11050 16510 11380
rect 16800 11050 16801 11380
rect 16509 11049 16801 11050
rect 17599 11380 17891 11381
rect 17599 11050 17600 11380
rect 17890 11050 17891 11380
rect 17599 11049 17891 11050
rect 18689 11380 18981 11381
rect 18689 11050 18690 11380
rect 18980 11050 18981 11380
rect 18689 11049 18981 11050
rect 19779 11380 20071 11381
rect 19779 11050 19780 11380
rect 20070 11050 20071 11380
rect 19779 11049 20071 11050
rect 20869 11380 21161 11381
rect 20869 11050 20870 11380
rect 21160 11050 21161 11380
rect 20869 11049 21161 11050
rect 179 11019 451 11020
rect 1240 2310 1450 2700
rect 5350 2321 5540 2920
rect 1240 2230 1250 2310
rect 1380 2230 1450 2310
rect 5349 2320 5541 2321
rect 1249 2229 1381 2230
rect 5349 2180 5350 2320
rect 5540 2180 5541 2320
rect 5349 2179 5541 2180
rect 379 450 761 451
rect 379 40 380 450
rect 760 40 761 450
rect 379 39 761 40
rect 1469 450 1851 451
rect 1469 40 1470 450
rect 1850 40 1851 450
rect 1469 39 1851 40
rect 2559 450 2941 451
rect 2559 40 2560 450
rect 2940 40 2941 450
rect 2559 39 2941 40
rect 3649 450 4031 451
rect 3649 40 3650 450
rect 4030 40 4031 450
rect 3649 39 4031 40
<< via4 >>
rect 180 11020 450 11390
rect 2330 11080 2620 11410
rect 3440 11080 3730 11410
rect 4490 11080 4780 11410
rect 5590 11080 5880 11410
rect 6700 11050 6990 11380
rect 7790 11050 8080 11380
rect 8880 11050 9170 11380
rect 9970 11050 10260 11380
rect 11060 11050 11350 11380
rect 12150 11050 12440 11380
rect 13240 11050 13530 11380
rect 14330 11050 14620 11380
rect 15420 11050 15710 11380
rect 16510 11050 16800 11380
rect 17600 11050 17890 11380
rect 18690 11050 18980 11380
rect 19780 11050 20070 11380
rect 20870 11050 21160 11380
rect 380 40 760 450
rect 1470 40 1850 450
rect 2560 40 2940 450
rect 3650 40 4030 450
<< metal5 >>
rect 2306 11430 2644 11434
rect 3416 11430 3754 11434
rect 4466 11430 4804 11434
rect 5566 11430 5904 11434
rect 150 11410 21770 11430
rect 150 11390 2330 11410
rect 150 11020 180 11390
rect 450 11080 2330 11390
rect 2620 11080 3440 11410
rect 3730 11080 4490 11410
rect 4780 11080 5590 11410
rect 5880 11380 21770 11410
rect 5880 11080 6700 11380
rect 450 11050 6700 11080
rect 6990 11050 7790 11380
rect 8080 11050 8880 11380
rect 9170 11050 9970 11380
rect 10260 11050 11060 11380
rect 11350 11050 12150 11380
rect 12440 11050 13240 11380
rect 13530 11050 14330 11380
rect 14620 11050 15420 11380
rect 15710 11050 16510 11380
rect 16800 11050 17600 11380
rect 17890 11050 18690 11380
rect 18980 11050 19780 11380
rect 20070 11050 20870 11380
rect 21160 11050 21770 11380
rect 450 11020 21770 11050
rect 150 10990 21770 11020
rect 3260 8710 3860 10990
rect 7250 8750 7850 10990
rect 11030 9970 11630 10990
rect 15090 10080 15690 10990
rect 10600 660 11320 3800
rect 14030 660 14750 3840
rect -20 450 19640 660
rect -20 40 380 450
rect 760 40 1470 450
rect 1850 40 2560 450
rect 2940 40 3650 450
rect 4030 40 19640 450
rect -20 10 19640 40
use bias_curm_n  bias_curm_n_0
timestamp 1654697490
transform 1 0 60 0 1 50
box -50 -50 1052 2198
use bias_curm_n  bias_curm_n_1
timestamp 1654697490
transform 1 0 1150 0 1 50
box -50 -50 1052 2198
use bias_curm_n  bias_curm_n_2
timestamp 1654697490
transform 1 0 2240 0 1 50
box -50 -50 1052 2198
use bias_curm_n  bias_curm_n_3
timestamp 1654697490
transform 1 0 3330 0 1 50
box -50 -50 1052 2198
use bias_curm_p  bias_curm_p_0
timestamp 1654704381
transform 1 0 20 0 1 3170
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_1
timestamp 1654704381
transform 1 0 1110 0 1 3170
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_2
timestamp 1654704381
transform 1 0 2200 0 1 3170
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_3
timestamp 1654704381
transform 1 0 2200 0 1 5460
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_4
timestamp 1654704381
transform 1 0 2200 0 1 7750
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_5
timestamp 1654704381
transform 1 0 2200 0 1 10040
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_6
timestamp 1654704381
transform 1 0 3290 0 1 10040
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_7
timestamp 1654704381
transform 1 0 20 0 1 5450
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_8
timestamp 1654704381
transform 1 0 5470 0 1 10040
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_9
timestamp 1654704381
transform 1 0 3290 0 1 7750
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_10
timestamp 1654704381
transform 1 0 3290 0 1 5460
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_11
timestamp 1654704381
transform 1 0 3290 0 1 3170
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_12
timestamp 1654704381
transform 1 0 5470 0 1 7750
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_13
timestamp 1654704381
transform 1 0 4380 0 1 7750
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_14
timestamp 1654704381
transform 1 0 4380 0 1 5460
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_15
timestamp 1654704381
transform 1 0 4380 0 1 3170
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_16
timestamp 1654704381
transform 1 0 5470 0 1 5460
box -10 -910 1100 1390
use bias_curm_p  bias_curm_p_17
timestamp 1654704381
transform 1 0 5470 0 1 3170
box -10 -910 1100 1390
use eight-mirrors-p  eight-mirrors-p_0
timestamp 1654704381
transform 1 0 6550 0 1 2260
box 0 0 2200 9140
use eight-mirrors-p  eight-mirrors-p_1
timestamp 1654704381
transform 1 0 8730 0 1 2260
box 0 0 2200 9140
use eight-mirrors-p  eight-mirrors-p_2
timestamp 1654704381
transform 1 0 13090 0 1 2260
box 0 0 2200 9140
use eight-mirrors-p  eight-mirrors-p_3
timestamp 1654704381
transform 1 0 10910 0 1 2260
box 0 0 2200 9140
use eight-mirrors-p  eight-mirrors-p_4
timestamp 1654704381
transform 1 0 17450 0 1 2260
box 0 0 2200 9140
use eight-mirrors-p  eight-mirrors-p_5
timestamp 1654704381
transform 1 0 15270 0 1 2260
box 0 0 2200 9140
use eight-mirrors-p  eight-mirrors-p_6
timestamp 1654704381
transform 1 0 19630 0 1 2260
box 0 0 2200 9140
use sky130_fd_pr__cap_mim_m3_2_26U9NK  sky130_fd_pr__cap_mim_m3_2_26U9NK_0
timestamp 1654701805
transform 0 1 2831 -1 0 5953
box -3351 -1601 3373 1601
use sky130_fd_pr__cap_mim_m3_2_26U9NK  sky130_fd_pr__cap_mim_m3_2_26U9NK_1
timestamp 1654701805
transform 0 1 6611 -1 0 5943
box -3351 -1601 3373 1601
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_1
timestamp 1654701805
transform 0 1 13261 -1 0 7053
box -3351 -3101 3373 3101
<< labels >>
rlabel metal5 4770 130 5030 460 1 VN
rlabel metal5 4960 11050 5220 11380 1 VP
rlabel metal3 40 2150 140 2250 1 I_in
rlabel metal3 670 5230 770 5330 1 FB_Bias_1
rlabel metal3 2860 2860 2980 3000 1 TIA_Bias
rlabel metal3 6150 2800 6290 2970 1 ctl_Bias
rlabel metal3 7570 2720 7750 2880 1 Comp_Bias_1
rlabel metal3 9730 2740 9880 2860 1 Comp_Bias_2
rlabel metal3 11910 2730 12060 2850 1 Comp_Bias_3
rlabel metal5 14070 2720 14220 2840 1 Comp_Bias_4
rlabel metal3 16330 2720 16470 2820 1 Comp_Bias_5
rlabel metal3 18470 2730 18610 2830 1 Comp_Bias_6
rlabel metal3 20660 2760 20840 2850 1 LVDS_Bias
rlabel metal3 4380 2800 4550 2940 1 Bias_Analog_out
rlabel metal4 5390 2330 5490 2420 1 vm12d
rlabel metal2 1040 2220 1130 2280 1 vm4d
<< end >>
