magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< metal3 >>
rect -3150 1072 3149 1100
rect -3150 -1072 3065 1072
rect 3129 -1072 3149 1072
rect -3150 -1100 3149 -1072
<< via3 >>
rect 3065 -1072 3129 1072
<< mimcap >>
rect -3050 960 2950 1000
rect -3050 -960 -3010 960
rect 2910 -960 2950 960
rect -3050 -1000 2950 -960
<< mimcapcontact >>
rect -3010 -960 2910 960
<< metal4 >>
rect 3049 1072 3145 1088
rect -3011 960 2911 961
rect -3011 -960 -3010 960
rect 2910 -960 2911 960
rect -3011 -961 2911 -960
rect 3049 -1072 3065 1072
rect 3129 -1072 3145 1072
rect 3049 -1088 3145 -1072
<< properties >>
string FIXED_BBOX -3150 -1100 3050 1100
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 10 val 615.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
