magic
tech sky130B
magscale 1 2
timestamp 1654633577
<< metal4 >>
rect -1351 1059 1351 1100
rect -1351 -1059 1095 1059
rect 1331 -1059 1351 1059
rect -1351 -1100 1351 -1059
<< via4 >>
rect 1095 -1059 1331 1059
<< mimcap2 >>
rect -1251 960 749 1000
rect -1251 -960 -1211 960
rect 709 -960 749 960
rect -1251 -1000 749 -960
<< mimcap2contact >>
rect -1211 -960 709 960
<< metal5 >>
rect 1053 1059 1373 1101
rect -1235 960 733 984
rect -1235 -960 -1211 960
rect 709 -960 733 960
rect -1235 -984 733 -960
rect 1053 -1059 1095 1059
rect 1331 -1059 1373 1059
rect 1053 -1101 1373 -1059
<< properties >>
string FIXED_BBOX -1351 -1100 849 1100
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10 l 10 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
