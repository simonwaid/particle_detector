magic
tech sky130A
magscale 1 2
timestamp 1647868710
<< error_p >>
rect -372 472 -314 478
rect -176 472 -118 478
rect 20 472 78 478
rect 216 472 274 478
rect 412 472 470 478
rect -372 438 -360 472
rect -176 438 -164 472
rect 20 438 32 472
rect 216 438 228 472
rect 412 438 424 472
rect -372 432 -314 438
rect -176 432 -118 438
rect 20 432 78 438
rect 216 432 274 438
rect 412 432 470 438
rect -470 -438 -412 -432
rect -274 -438 -216 -432
rect -78 -438 -20 -432
rect 118 -438 176 -432
rect 314 -438 372 -432
rect -470 -472 -458 -438
rect -274 -472 -262 -438
rect -78 -472 -66 -438
rect 118 -472 130 -438
rect 314 -472 326 -438
rect -470 -478 -412 -472
rect -274 -478 -216 -472
rect -78 -478 -20 -472
rect 118 -478 176 -472
rect 314 -478 372 -472
<< pwell >>
rect -657 -610 657 610
<< nmoslvt >>
rect -461 -400 -421 400
rect -363 -400 -323 400
rect -265 -400 -225 400
rect -167 -400 -127 400
rect -69 -400 -29 400
rect 29 -400 69 400
rect 127 -400 167 400
rect 225 -400 265 400
rect 323 -400 363 400
rect 421 -400 461 400
<< ndiff >>
rect -519 388 -461 400
rect -519 -388 -507 388
rect -473 -388 -461 388
rect -519 -400 -461 -388
rect -421 388 -363 400
rect -421 -388 -409 388
rect -375 -388 -363 388
rect -421 -400 -363 -388
rect -323 388 -265 400
rect -323 -388 -311 388
rect -277 -388 -265 388
rect -323 -400 -265 -388
rect -225 388 -167 400
rect -225 -388 -213 388
rect -179 -388 -167 388
rect -225 -400 -167 -388
rect -127 388 -69 400
rect -127 -388 -115 388
rect -81 -388 -69 388
rect -127 -400 -69 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 69 388 127 400
rect 69 -388 81 388
rect 115 -388 127 388
rect 69 -400 127 -388
rect 167 388 225 400
rect 167 -388 179 388
rect 213 -388 225 388
rect 167 -400 225 -388
rect 265 388 323 400
rect 265 -388 277 388
rect 311 -388 323 388
rect 265 -400 323 -388
rect 363 388 421 400
rect 363 -388 375 388
rect 409 -388 421 388
rect 363 -400 421 -388
rect 461 388 519 400
rect 461 -388 473 388
rect 507 -388 519 388
rect 461 -400 519 -388
<< ndiffc >>
rect -507 -388 -473 388
rect -409 -388 -375 388
rect -311 -388 -277 388
rect -213 -388 -179 388
rect -115 -388 -81 388
rect -17 -388 17 388
rect 81 -388 115 388
rect 179 -388 213 388
rect 277 -388 311 388
rect 375 -388 409 388
rect 473 -388 507 388
<< psubdiff >>
rect -621 540 -525 574
rect 525 540 621 574
rect -621 478 -587 540
rect 587 478 621 540
rect -621 -540 -587 -478
rect 587 -540 621 -478
rect -621 -574 -525 -540
rect 525 -574 621 -540
<< psubdiffcont >>
rect -525 540 525 574
rect -621 -478 -587 478
rect 587 -478 621 478
rect -525 -574 525 -540
<< poly >>
rect -376 472 -310 488
rect -376 438 -360 472
rect -326 438 -310 472
rect -461 400 -421 426
rect -376 422 -310 438
rect -180 472 -114 488
rect -180 438 -164 472
rect -130 438 -114 472
rect -363 400 -323 422
rect -265 400 -225 426
rect -180 422 -114 438
rect 16 472 82 488
rect 16 438 32 472
rect 66 438 82 472
rect -167 400 -127 422
rect -69 400 -29 426
rect 16 422 82 438
rect 212 472 278 488
rect 212 438 228 472
rect 262 438 278 472
rect 29 400 69 422
rect 127 400 167 426
rect 212 422 278 438
rect 408 472 474 488
rect 408 438 424 472
rect 458 438 474 472
rect 225 400 265 422
rect 323 400 363 426
rect 408 422 474 438
rect 421 400 461 422
rect -461 -422 -421 -400
rect -474 -438 -408 -422
rect -363 -426 -323 -400
rect -265 -422 -225 -400
rect -474 -472 -458 -438
rect -424 -472 -408 -438
rect -474 -488 -408 -472
rect -278 -438 -212 -422
rect -167 -426 -127 -400
rect -69 -422 -29 -400
rect -278 -472 -262 -438
rect -228 -472 -212 -438
rect -278 -488 -212 -472
rect -82 -438 -16 -422
rect 29 -426 69 -400
rect 127 -422 167 -400
rect -82 -472 -66 -438
rect -32 -472 -16 -438
rect -82 -488 -16 -472
rect 114 -438 180 -422
rect 225 -426 265 -400
rect 323 -422 363 -400
rect 114 -472 130 -438
rect 164 -472 180 -438
rect 114 -488 180 -472
rect 310 -438 376 -422
rect 421 -426 461 -400
rect 310 -472 326 -438
rect 360 -472 376 -438
rect 310 -488 376 -472
<< polycont >>
rect -360 438 -326 472
rect -164 438 -130 472
rect 32 438 66 472
rect 228 438 262 472
rect 424 438 458 472
rect -458 -472 -424 -438
rect -262 -472 -228 -438
rect -66 -472 -32 -438
rect 130 -472 164 -438
rect 326 -472 360 -438
<< locali >>
rect -621 540 -525 574
rect 525 540 621 574
rect -621 478 -587 540
rect 587 478 621 540
rect -376 438 -360 472
rect -326 438 -310 472
rect -180 438 -164 472
rect -130 438 -114 472
rect 16 438 32 472
rect 66 438 82 472
rect 212 438 228 472
rect 262 438 278 472
rect 408 438 424 472
rect 458 438 474 472
rect -507 388 -473 404
rect -507 -404 -473 -388
rect -409 388 -375 404
rect -409 -404 -375 -388
rect -311 388 -277 404
rect -311 -404 -277 -388
rect -213 388 -179 404
rect -213 -404 -179 -388
rect -115 388 -81 404
rect -115 -404 -81 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 81 388 115 404
rect 81 -404 115 -388
rect 179 388 213 404
rect 179 -404 213 -388
rect 277 388 311 404
rect 277 -404 311 -388
rect 375 388 409 404
rect 375 -404 409 -388
rect 473 388 507 404
rect 473 -404 507 -388
rect -474 -472 -458 -438
rect -424 -472 -408 -438
rect -278 -472 -262 -438
rect -228 -472 -212 -438
rect -82 -472 -66 -438
rect -32 -472 -16 -438
rect 114 -472 130 -438
rect 164 -472 180 -438
rect 310 -472 326 -438
rect 360 -472 376 -438
rect -621 -540 -587 -478
rect 587 -540 621 -478
rect -621 -574 -525 -540
rect 525 -574 621 -540
<< viali >>
rect -360 438 -326 472
rect -164 438 -130 472
rect 32 438 66 472
rect 228 438 262 472
rect 424 438 458 472
rect -507 -388 -473 388
rect -409 -388 -375 388
rect -311 -388 -277 388
rect -213 -388 -179 388
rect -115 -388 -81 388
rect -17 -388 17 388
rect 81 -388 115 388
rect 179 -388 213 388
rect 277 -388 311 388
rect 375 -388 409 388
rect 473 -388 507 388
rect -458 -472 -424 -438
rect -262 -472 -228 -438
rect -66 -472 -32 -438
rect 130 -472 164 -438
rect 326 -472 360 -438
<< metal1 >>
rect -372 472 -314 478
rect -372 438 -360 472
rect -326 438 -314 472
rect -372 432 -314 438
rect -176 472 -118 478
rect -176 438 -164 472
rect -130 438 -118 472
rect -176 432 -118 438
rect 20 472 78 478
rect 20 438 32 472
rect 66 438 78 472
rect 20 432 78 438
rect 216 472 274 478
rect 216 438 228 472
rect 262 438 274 472
rect 216 432 274 438
rect 412 472 470 478
rect 412 438 424 472
rect 458 438 470 472
rect 412 432 470 438
rect -513 388 -467 400
rect -513 -388 -507 388
rect -473 -388 -467 388
rect -513 -400 -467 -388
rect -415 388 -369 400
rect -415 -388 -409 388
rect -375 -388 -369 388
rect -415 -400 -369 -388
rect -317 388 -271 400
rect -317 -388 -311 388
rect -277 -388 -271 388
rect -317 -400 -271 -388
rect -219 388 -173 400
rect -219 -388 -213 388
rect -179 -388 -173 388
rect -219 -400 -173 -388
rect -121 388 -75 400
rect -121 -388 -115 388
rect -81 -388 -75 388
rect -121 -400 -75 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 75 388 121 400
rect 75 -388 81 388
rect 115 -388 121 388
rect 75 -400 121 -388
rect 173 388 219 400
rect 173 -388 179 388
rect 213 -388 219 388
rect 173 -400 219 -388
rect 271 388 317 400
rect 271 -388 277 388
rect 311 -388 317 388
rect 271 -400 317 -388
rect 369 388 415 400
rect 369 -388 375 388
rect 409 -388 415 388
rect 369 -400 415 -388
rect 467 388 513 400
rect 467 -388 473 388
rect 507 -388 513 388
rect 467 -400 513 -388
rect -470 -438 -412 -432
rect -470 -472 -458 -438
rect -424 -472 -412 -438
rect -470 -478 -412 -472
rect -274 -438 -216 -432
rect -274 -472 -262 -438
rect -228 -472 -216 -438
rect -274 -478 -216 -472
rect -78 -438 -20 -432
rect -78 -472 -66 -438
rect -32 -472 -20 -438
rect -78 -478 -20 -472
rect 118 -438 176 -432
rect 118 -472 130 -438
rect 164 -472 176 -438
rect 118 -478 176 -472
rect 314 -438 372 -432
rect 314 -472 326 -438
rect 360 -472 372 -438
rect 314 -478 372 -472
<< properties >>
string FIXED_BBOX -604 -557 604 557
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4 l 0.2 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
