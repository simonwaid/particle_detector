magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< nwell >>
rect -957 -419 957 419
<< pmos >>
rect -761 -200 -661 200
rect -603 -200 -503 200
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
rect 503 -200 603 200
rect 661 -200 761 200
<< pdiff >>
rect -819 188 -761 200
rect -819 -188 -807 188
rect -773 -188 -761 188
rect -819 -200 -761 -188
rect -661 188 -603 200
rect -661 -188 -649 188
rect -615 -188 -603 188
rect -661 -200 -603 -188
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
rect 603 188 661 200
rect 603 -188 615 188
rect 649 -188 661 188
rect 603 -200 661 -188
rect 761 188 819 200
rect 761 -188 773 188
rect 807 -188 819 188
rect 761 -200 819 -188
<< pdiffc >>
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
<< nsubdiff >>
rect -921 349 -825 383
rect 825 349 921 383
rect -921 287 -887 349
rect 887 287 921 349
rect -921 -349 -887 -287
rect 887 -349 921 -287
rect -921 -383 -825 -349
rect 825 -383 921 -349
<< nsubdiffcont >>
rect -825 349 825 383
rect -921 -287 -887 287
rect 887 -287 921 287
rect -825 -383 825 -349
<< poly >>
rect -761 281 -661 297
rect -761 247 -745 281
rect -677 247 -661 281
rect -761 200 -661 247
rect -603 281 -503 297
rect -603 247 -587 281
rect -519 247 -503 281
rect -603 200 -503 247
rect -445 281 -345 297
rect -445 247 -429 281
rect -361 247 -345 281
rect -445 200 -345 247
rect -287 281 -187 297
rect -287 247 -271 281
rect -203 247 -187 281
rect -287 200 -187 247
rect -129 281 -29 297
rect -129 247 -113 281
rect -45 247 -29 281
rect -129 200 -29 247
rect 29 281 129 297
rect 29 247 45 281
rect 113 247 129 281
rect 29 200 129 247
rect 187 281 287 297
rect 187 247 203 281
rect 271 247 287 281
rect 187 200 287 247
rect 345 281 445 297
rect 345 247 361 281
rect 429 247 445 281
rect 345 200 445 247
rect 503 281 603 297
rect 503 247 519 281
rect 587 247 603 281
rect 503 200 603 247
rect 661 281 761 297
rect 661 247 677 281
rect 745 247 761 281
rect 661 200 761 247
rect -761 -247 -661 -200
rect -761 -281 -745 -247
rect -677 -281 -661 -247
rect -761 -297 -661 -281
rect -603 -247 -503 -200
rect -603 -281 -587 -247
rect -519 -281 -503 -247
rect -603 -297 -503 -281
rect -445 -247 -345 -200
rect -445 -281 -429 -247
rect -361 -281 -345 -247
rect -445 -297 -345 -281
rect -287 -247 -187 -200
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -287 -297 -187 -281
rect -129 -247 -29 -200
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect -129 -297 -29 -281
rect 29 -247 129 -200
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 29 -297 129 -281
rect 187 -247 287 -200
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 187 -297 287 -281
rect 345 -247 445 -200
rect 345 -281 361 -247
rect 429 -281 445 -247
rect 345 -297 445 -281
rect 503 -247 603 -200
rect 503 -281 519 -247
rect 587 -281 603 -247
rect 503 -297 603 -281
rect 661 -247 761 -200
rect 661 -281 677 -247
rect 745 -281 761 -247
rect 661 -297 761 -281
<< polycont >>
rect -745 247 -677 281
rect -587 247 -519 281
rect -429 247 -361 281
rect -271 247 -203 281
rect -113 247 -45 281
rect 45 247 113 281
rect 203 247 271 281
rect 361 247 429 281
rect 519 247 587 281
rect 677 247 745 281
rect -745 -281 -677 -247
rect -587 -281 -519 -247
rect -429 -281 -361 -247
rect -271 -281 -203 -247
rect -113 -281 -45 -247
rect 45 -281 113 -247
rect 203 -281 271 -247
rect 361 -281 429 -247
rect 519 -281 587 -247
rect 677 -281 745 -247
<< locali >>
rect -921 349 -825 383
rect 825 349 921 383
rect -921 287 -887 349
rect 887 287 921 349
rect -761 247 -745 281
rect -677 247 -661 281
rect -603 247 -587 281
rect -519 247 -503 281
rect -445 247 -429 281
rect -361 247 -345 281
rect -287 247 -271 281
rect -203 247 -187 281
rect -129 247 -113 281
rect -45 247 -29 281
rect 29 247 45 281
rect 113 247 129 281
rect 187 247 203 281
rect 271 247 287 281
rect 345 247 361 281
rect 429 247 445 281
rect 503 247 519 281
rect 587 247 603 281
rect 661 247 677 281
rect 745 247 761 281
rect -807 188 -773 204
rect -807 -204 -773 -188
rect -649 188 -615 204
rect -649 -204 -615 -188
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect 615 188 649 204
rect 615 -204 649 -188
rect 773 188 807 204
rect 773 -204 807 -188
rect -761 -281 -745 -247
rect -677 -281 -661 -247
rect -603 -281 -587 -247
rect -519 -281 -503 -247
rect -445 -281 -429 -247
rect -361 -281 -345 -247
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 345 -281 361 -247
rect 429 -281 445 -247
rect 503 -281 519 -247
rect 587 -281 603 -247
rect 661 -281 677 -247
rect 745 -281 761 -247
rect -921 -349 -887 -287
rect 887 -349 921 -287
rect -921 -383 -825 -349
rect 825 -383 921 -349
<< viali >>
rect -745 247 -677 281
rect -587 247 -519 281
rect -429 247 -361 281
rect -271 247 -203 281
rect -113 247 -45 281
rect 45 247 113 281
rect 203 247 271 281
rect 361 247 429 281
rect 519 247 587 281
rect 677 247 745 281
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect -745 -281 -677 -247
rect -587 -281 -519 -247
rect -429 -281 -361 -247
rect -271 -281 -203 -247
rect -113 -281 -45 -247
rect 45 -281 113 -247
rect 203 -281 271 -247
rect 361 -281 429 -247
rect 519 -281 587 -247
rect 677 -281 745 -247
<< metal1 >>
rect -757 281 -665 287
rect -757 247 -745 281
rect -677 247 -665 281
rect -757 241 -665 247
rect -599 281 -507 287
rect -599 247 -587 281
rect -519 247 -507 281
rect -599 241 -507 247
rect -441 281 -349 287
rect -441 247 -429 281
rect -361 247 -349 281
rect -441 241 -349 247
rect -283 281 -191 287
rect -283 247 -271 281
rect -203 247 -191 281
rect -283 241 -191 247
rect -125 281 -33 287
rect -125 247 -113 281
rect -45 247 -33 281
rect -125 241 -33 247
rect 33 281 125 287
rect 33 247 45 281
rect 113 247 125 281
rect 33 241 125 247
rect 191 281 283 287
rect 191 247 203 281
rect 271 247 283 281
rect 191 241 283 247
rect 349 281 441 287
rect 349 247 361 281
rect 429 247 441 281
rect 349 241 441 247
rect 507 281 599 287
rect 507 247 519 281
rect 587 247 599 281
rect 507 241 599 247
rect 665 281 757 287
rect 665 247 677 281
rect 745 247 757 281
rect 665 241 757 247
rect -813 188 -767 200
rect -813 -188 -807 188
rect -773 -188 -767 188
rect -813 -200 -767 -188
rect -655 188 -609 200
rect -655 -188 -649 188
rect -615 -188 -609 188
rect -655 -200 -609 -188
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect 609 188 655 200
rect 609 -188 615 188
rect 649 -188 655 188
rect 609 -200 655 -188
rect 767 188 813 200
rect 767 -188 773 188
rect 807 -188 813 188
rect 767 -200 813 -188
rect -757 -247 -665 -241
rect -757 -281 -745 -247
rect -677 -281 -665 -247
rect -757 -287 -665 -281
rect -599 -247 -507 -241
rect -599 -281 -587 -247
rect -519 -281 -507 -247
rect -599 -287 -507 -281
rect -441 -247 -349 -241
rect -441 -281 -429 -247
rect -361 -281 -349 -247
rect -441 -287 -349 -281
rect -283 -247 -191 -241
rect -283 -281 -271 -247
rect -203 -281 -191 -247
rect -283 -287 -191 -281
rect -125 -247 -33 -241
rect -125 -281 -113 -247
rect -45 -281 -33 -247
rect -125 -287 -33 -281
rect 33 -247 125 -241
rect 33 -281 45 -247
rect 113 -281 125 -247
rect 33 -287 125 -281
rect 191 -247 283 -241
rect 191 -281 203 -247
rect 271 -281 283 -247
rect 191 -287 283 -281
rect 349 -247 441 -241
rect 349 -281 361 -247
rect 429 -281 441 -247
rect 349 -287 441 -281
rect 507 -247 599 -241
rect 507 -281 519 -247
rect 587 -281 599 -247
rect 507 -287 599 -281
rect 665 -247 757 -241
rect 665 -281 677 -247
rect 745 -281 757 -247
rect 665 -287 757 -281
<< properties >>
string FIXED_BBOX -904 -366 904 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
