magic
tech sky130A
magscale 1 2
timestamp 1645802395
<< metal4 >>
rect -3351 659 3351 700
rect -3351 -659 3095 659
rect 3331 -659 3351 659
rect -3351 -700 3351 -659
<< via4 >>
rect 3095 -659 3331 659
<< mimcap2 >>
rect -3251 560 2749 600
rect -3251 -560 -3211 560
rect 2709 -560 2749 560
rect -3251 -600 2749 -560
<< mimcap2contact >>
rect -3211 -560 2709 560
<< metal5 >>
rect 3053 659 3373 701
rect -3235 560 2733 584
rect -3235 -560 -3211 560
rect 2709 -560 2733 560
rect -3235 -584 2733 -560
rect 3053 -659 3095 659
rect 3331 -659 3373 659
rect 3053 -701 3373 -659
<< properties >>
string FIXED_BBOX -3351 -700 2849 700
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 6 val 373.68 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
