magic
tech sky130A
timestamp 1647868710
<< metal2 >>
rect 5935 5190 7170 5275
rect 13075 5190 14310 5275
rect 20200 5190 21435 5275
rect 5955 4555 7190 4640
rect 13075 4555 14310 4640
rect 20200 4555 21435 4640
rect 6490 4080 7220 4160
rect 13620 4080 14350 4160
rect 20745 4080 21475 4160
<< metal3 >>
rect 5845 7120 27355 7490
rect 1040 4245 1140 4310
rect 6505 4205 7685 4275
rect 6505 4200 7110 4205
rect 7605 4200 7685 4205
rect 13605 4205 14795 4280
rect 13605 4195 14265 4205
rect 14725 4195 14795 4205
rect 20740 4210 21930 4285
rect 20740 4200 21390 4210
rect 21850 4200 21930 4210
rect 7080 -10 7155 500
rect 14205 -10 14280 500
rect 21330 -10 21405 500
<< metal4 >>
rect 5985 6440 7840 6720
rect 13110 6440 14885 6720
rect 20235 6440 22010 6720
rect 5985 6100 7840 6380
rect 13110 6100 14885 6380
rect 20235 6100 22010 6380
use outd_stage2  outd_stage2_0
timestamp 1647868710
transform 1 0 5 0 1 430
box -15 -440 7116 7060
use outd_stage2  outd_stage2_1
timestamp 1647868710
transform 1 0 7130 0 1 430
box -15 -440 7116 7060
use outd_stage2  outd_stage2_2
timestamp 1647868710
transform 1 0 14255 0 1 430
box -15 -440 7116 7060
use outd_stage2  outd_stage2_3
timestamp 1647868710
transform 1 0 21380 0 1 430
box -15 -440 7116 7060
<< end >>
