magic
tech sky130A
magscale 1 2
timestamp 1645790779
<< error_p >>
rect -2381 581 -2323 587
rect -2189 581 -2131 587
rect -1997 581 -1939 587
rect -1805 581 -1747 587
rect -1613 581 -1555 587
rect -1421 581 -1363 587
rect -1229 581 -1171 587
rect -1037 581 -979 587
rect -845 581 -787 587
rect -653 581 -595 587
rect -461 581 -403 587
rect -269 581 -211 587
rect -77 581 -19 587
rect 115 581 173 587
rect 307 581 365 587
rect 499 581 557 587
rect 691 581 749 587
rect 883 581 941 587
rect 1075 581 1133 587
rect 1267 581 1325 587
rect 1459 581 1517 587
rect 1651 581 1709 587
rect 1843 581 1901 587
rect 2035 581 2093 587
rect 2227 581 2285 587
rect -2381 547 -2369 581
rect -2189 547 -2177 581
rect -1997 547 -1985 581
rect -1805 547 -1793 581
rect -1613 547 -1601 581
rect -1421 547 -1409 581
rect -1229 547 -1217 581
rect -1037 547 -1025 581
rect -845 547 -833 581
rect -653 547 -641 581
rect -461 547 -449 581
rect -269 547 -257 581
rect -77 547 -65 581
rect 115 547 127 581
rect 307 547 319 581
rect 499 547 511 581
rect 691 547 703 581
rect 883 547 895 581
rect 1075 547 1087 581
rect 1267 547 1279 581
rect 1459 547 1471 581
rect 1651 547 1663 581
rect 1843 547 1855 581
rect 2035 547 2047 581
rect 2227 547 2239 581
rect -2381 541 -2323 547
rect -2189 541 -2131 547
rect -1997 541 -1939 547
rect -1805 541 -1747 547
rect -1613 541 -1555 547
rect -1421 541 -1363 547
rect -1229 541 -1171 547
rect -1037 541 -979 547
rect -845 541 -787 547
rect -653 541 -595 547
rect -461 541 -403 547
rect -269 541 -211 547
rect -77 541 -19 547
rect 115 541 173 547
rect 307 541 365 547
rect 499 541 557 547
rect 691 541 749 547
rect 883 541 941 547
rect 1075 541 1133 547
rect 1267 541 1325 547
rect 1459 541 1517 547
rect 1651 541 1709 547
rect 1843 541 1901 547
rect 2035 541 2093 547
rect 2227 541 2285 547
rect -2285 71 -2227 77
rect -2093 71 -2035 77
rect -1901 71 -1843 77
rect -1709 71 -1651 77
rect -1517 71 -1459 77
rect -1325 71 -1267 77
rect -1133 71 -1075 77
rect -941 71 -883 77
rect -749 71 -691 77
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect 595 71 653 77
rect 787 71 845 77
rect 979 71 1037 77
rect 1171 71 1229 77
rect 1363 71 1421 77
rect 1555 71 1613 77
rect 1747 71 1805 77
rect 1939 71 1997 77
rect 2131 71 2189 77
rect 2323 71 2381 77
rect -2285 37 -2273 71
rect -2093 37 -2081 71
rect -1901 37 -1889 71
rect -1709 37 -1697 71
rect -1517 37 -1505 71
rect -1325 37 -1313 71
rect -1133 37 -1121 71
rect -941 37 -929 71
rect -749 37 -737 71
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect 595 37 607 71
rect 787 37 799 71
rect 979 37 991 71
rect 1171 37 1183 71
rect 1363 37 1375 71
rect 1555 37 1567 71
rect 1747 37 1759 71
rect 1939 37 1951 71
rect 2131 37 2143 71
rect 2323 37 2335 71
rect -2285 31 -2227 37
rect -2093 31 -2035 37
rect -1901 31 -1843 37
rect -1709 31 -1651 37
rect -1517 31 -1459 37
rect -1325 31 -1267 37
rect -1133 31 -1075 37
rect -941 31 -883 37
rect -749 31 -691 37
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect 595 31 653 37
rect 787 31 845 37
rect 979 31 1037 37
rect 1171 31 1229 37
rect 1363 31 1421 37
rect 1555 31 1613 37
rect 1747 31 1805 37
rect 1939 31 1997 37
rect 2131 31 2189 37
rect 2323 31 2381 37
rect -2285 -37 -2227 -31
rect -2093 -37 -2035 -31
rect -1901 -37 -1843 -31
rect -1709 -37 -1651 -31
rect -1517 -37 -1459 -31
rect -1325 -37 -1267 -31
rect -1133 -37 -1075 -31
rect -941 -37 -883 -31
rect -749 -37 -691 -31
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect 595 -37 653 -31
rect 787 -37 845 -31
rect 979 -37 1037 -31
rect 1171 -37 1229 -31
rect 1363 -37 1421 -31
rect 1555 -37 1613 -31
rect 1747 -37 1805 -31
rect 1939 -37 1997 -31
rect 2131 -37 2189 -31
rect 2323 -37 2381 -31
rect -2285 -71 -2273 -37
rect -2093 -71 -2081 -37
rect -1901 -71 -1889 -37
rect -1709 -71 -1697 -37
rect -1517 -71 -1505 -37
rect -1325 -71 -1313 -37
rect -1133 -71 -1121 -37
rect -941 -71 -929 -37
rect -749 -71 -737 -37
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect 595 -71 607 -37
rect 787 -71 799 -37
rect 979 -71 991 -37
rect 1171 -71 1183 -37
rect 1363 -71 1375 -37
rect 1555 -71 1567 -37
rect 1747 -71 1759 -37
rect 1939 -71 1951 -37
rect 2131 -71 2143 -37
rect 2323 -71 2335 -37
rect -2285 -77 -2227 -71
rect -2093 -77 -2035 -71
rect -1901 -77 -1843 -71
rect -1709 -77 -1651 -71
rect -1517 -77 -1459 -71
rect -1325 -77 -1267 -71
rect -1133 -77 -1075 -71
rect -941 -77 -883 -71
rect -749 -77 -691 -71
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect 595 -77 653 -71
rect 787 -77 845 -71
rect 979 -77 1037 -71
rect 1171 -77 1229 -71
rect 1363 -77 1421 -71
rect 1555 -77 1613 -71
rect 1747 -77 1805 -71
rect 1939 -77 1997 -71
rect 2131 -77 2189 -71
rect 2323 -77 2381 -71
rect -2381 -547 -2323 -541
rect -2189 -547 -2131 -541
rect -1997 -547 -1939 -541
rect -1805 -547 -1747 -541
rect -1613 -547 -1555 -541
rect -1421 -547 -1363 -541
rect -1229 -547 -1171 -541
rect -1037 -547 -979 -541
rect -845 -547 -787 -541
rect -653 -547 -595 -541
rect -461 -547 -403 -541
rect -269 -547 -211 -541
rect -77 -547 -19 -541
rect 115 -547 173 -541
rect 307 -547 365 -541
rect 499 -547 557 -541
rect 691 -547 749 -541
rect 883 -547 941 -541
rect 1075 -547 1133 -541
rect 1267 -547 1325 -541
rect 1459 -547 1517 -541
rect 1651 -547 1709 -541
rect 1843 -547 1901 -541
rect 2035 -547 2093 -541
rect 2227 -547 2285 -541
rect -2381 -581 -2369 -547
rect -2189 -581 -2177 -547
rect -1997 -581 -1985 -547
rect -1805 -581 -1793 -547
rect -1613 -581 -1601 -547
rect -1421 -581 -1409 -547
rect -1229 -581 -1217 -547
rect -1037 -581 -1025 -547
rect -845 -581 -833 -547
rect -653 -581 -641 -547
rect -461 -581 -449 -547
rect -269 -581 -257 -547
rect -77 -581 -65 -547
rect 115 -581 127 -547
rect 307 -581 319 -547
rect 499 -581 511 -547
rect 691 -581 703 -547
rect 883 -581 895 -547
rect 1075 -581 1087 -547
rect 1267 -581 1279 -547
rect 1459 -581 1471 -547
rect 1651 -581 1663 -547
rect 1843 -581 1855 -547
rect 2035 -581 2047 -547
rect 2227 -581 2239 -547
rect -2381 -587 -2323 -581
rect -2189 -587 -2131 -581
rect -1997 -587 -1939 -581
rect -1805 -587 -1747 -581
rect -1613 -587 -1555 -581
rect -1421 -587 -1363 -581
rect -1229 -587 -1171 -581
rect -1037 -587 -979 -581
rect -845 -587 -787 -581
rect -653 -587 -595 -581
rect -461 -587 -403 -581
rect -269 -587 -211 -581
rect -77 -587 -19 -581
rect 115 -587 173 -581
rect 307 -587 365 -581
rect 499 -587 557 -581
rect 691 -587 749 -581
rect 883 -587 941 -581
rect 1075 -587 1133 -581
rect 1267 -587 1325 -581
rect 1459 -587 1517 -581
rect 1651 -587 1709 -581
rect 1843 -587 1901 -581
rect 2035 -587 2093 -581
rect 2227 -587 2285 -581
<< pwell >>
rect -2567 -719 2567 719
<< nmos >>
rect -2367 109 -2337 509
rect -2271 109 -2241 509
rect -2175 109 -2145 509
rect -2079 109 -2049 509
rect -1983 109 -1953 509
rect -1887 109 -1857 509
rect -1791 109 -1761 509
rect -1695 109 -1665 509
rect -1599 109 -1569 509
rect -1503 109 -1473 509
rect -1407 109 -1377 509
rect -1311 109 -1281 509
rect -1215 109 -1185 509
rect -1119 109 -1089 509
rect -1023 109 -993 509
rect -927 109 -897 509
rect -831 109 -801 509
rect -735 109 -705 509
rect -639 109 -609 509
rect -543 109 -513 509
rect -447 109 -417 509
rect -351 109 -321 509
rect -255 109 -225 509
rect -159 109 -129 509
rect -63 109 -33 509
rect 33 109 63 509
rect 129 109 159 509
rect 225 109 255 509
rect 321 109 351 509
rect 417 109 447 509
rect 513 109 543 509
rect 609 109 639 509
rect 705 109 735 509
rect 801 109 831 509
rect 897 109 927 509
rect 993 109 1023 509
rect 1089 109 1119 509
rect 1185 109 1215 509
rect 1281 109 1311 509
rect 1377 109 1407 509
rect 1473 109 1503 509
rect 1569 109 1599 509
rect 1665 109 1695 509
rect 1761 109 1791 509
rect 1857 109 1887 509
rect 1953 109 1983 509
rect 2049 109 2079 509
rect 2145 109 2175 509
rect 2241 109 2271 509
rect 2337 109 2367 509
rect -2367 -509 -2337 -109
rect -2271 -509 -2241 -109
rect -2175 -509 -2145 -109
rect -2079 -509 -2049 -109
rect -1983 -509 -1953 -109
rect -1887 -509 -1857 -109
rect -1791 -509 -1761 -109
rect -1695 -509 -1665 -109
rect -1599 -509 -1569 -109
rect -1503 -509 -1473 -109
rect -1407 -509 -1377 -109
rect -1311 -509 -1281 -109
rect -1215 -509 -1185 -109
rect -1119 -509 -1089 -109
rect -1023 -509 -993 -109
rect -927 -509 -897 -109
rect -831 -509 -801 -109
rect -735 -509 -705 -109
rect -639 -509 -609 -109
rect -543 -509 -513 -109
rect -447 -509 -417 -109
rect -351 -509 -321 -109
rect -255 -509 -225 -109
rect -159 -509 -129 -109
rect -63 -509 -33 -109
rect 33 -509 63 -109
rect 129 -509 159 -109
rect 225 -509 255 -109
rect 321 -509 351 -109
rect 417 -509 447 -109
rect 513 -509 543 -109
rect 609 -509 639 -109
rect 705 -509 735 -109
rect 801 -509 831 -109
rect 897 -509 927 -109
rect 993 -509 1023 -109
rect 1089 -509 1119 -109
rect 1185 -509 1215 -109
rect 1281 -509 1311 -109
rect 1377 -509 1407 -109
rect 1473 -509 1503 -109
rect 1569 -509 1599 -109
rect 1665 -509 1695 -109
rect 1761 -509 1791 -109
rect 1857 -509 1887 -109
rect 1953 -509 1983 -109
rect 2049 -509 2079 -109
rect 2145 -509 2175 -109
rect 2241 -509 2271 -109
rect 2337 -509 2367 -109
<< ndiff >>
rect -2429 497 -2367 509
rect -2429 121 -2417 497
rect -2383 121 -2367 497
rect -2429 109 -2367 121
rect -2337 497 -2271 509
rect -2337 121 -2321 497
rect -2287 121 -2271 497
rect -2337 109 -2271 121
rect -2241 497 -2175 509
rect -2241 121 -2225 497
rect -2191 121 -2175 497
rect -2241 109 -2175 121
rect -2145 497 -2079 509
rect -2145 121 -2129 497
rect -2095 121 -2079 497
rect -2145 109 -2079 121
rect -2049 497 -1983 509
rect -2049 121 -2033 497
rect -1999 121 -1983 497
rect -2049 109 -1983 121
rect -1953 497 -1887 509
rect -1953 121 -1937 497
rect -1903 121 -1887 497
rect -1953 109 -1887 121
rect -1857 497 -1791 509
rect -1857 121 -1841 497
rect -1807 121 -1791 497
rect -1857 109 -1791 121
rect -1761 497 -1695 509
rect -1761 121 -1745 497
rect -1711 121 -1695 497
rect -1761 109 -1695 121
rect -1665 497 -1599 509
rect -1665 121 -1649 497
rect -1615 121 -1599 497
rect -1665 109 -1599 121
rect -1569 497 -1503 509
rect -1569 121 -1553 497
rect -1519 121 -1503 497
rect -1569 109 -1503 121
rect -1473 497 -1407 509
rect -1473 121 -1457 497
rect -1423 121 -1407 497
rect -1473 109 -1407 121
rect -1377 497 -1311 509
rect -1377 121 -1361 497
rect -1327 121 -1311 497
rect -1377 109 -1311 121
rect -1281 497 -1215 509
rect -1281 121 -1265 497
rect -1231 121 -1215 497
rect -1281 109 -1215 121
rect -1185 497 -1119 509
rect -1185 121 -1169 497
rect -1135 121 -1119 497
rect -1185 109 -1119 121
rect -1089 497 -1023 509
rect -1089 121 -1073 497
rect -1039 121 -1023 497
rect -1089 109 -1023 121
rect -993 497 -927 509
rect -993 121 -977 497
rect -943 121 -927 497
rect -993 109 -927 121
rect -897 497 -831 509
rect -897 121 -881 497
rect -847 121 -831 497
rect -897 109 -831 121
rect -801 497 -735 509
rect -801 121 -785 497
rect -751 121 -735 497
rect -801 109 -735 121
rect -705 497 -639 509
rect -705 121 -689 497
rect -655 121 -639 497
rect -705 109 -639 121
rect -609 497 -543 509
rect -609 121 -593 497
rect -559 121 -543 497
rect -609 109 -543 121
rect -513 497 -447 509
rect -513 121 -497 497
rect -463 121 -447 497
rect -513 109 -447 121
rect -417 497 -351 509
rect -417 121 -401 497
rect -367 121 -351 497
rect -417 109 -351 121
rect -321 497 -255 509
rect -321 121 -305 497
rect -271 121 -255 497
rect -321 109 -255 121
rect -225 497 -159 509
rect -225 121 -209 497
rect -175 121 -159 497
rect -225 109 -159 121
rect -129 497 -63 509
rect -129 121 -113 497
rect -79 121 -63 497
rect -129 109 -63 121
rect -33 497 33 509
rect -33 121 -17 497
rect 17 121 33 497
rect -33 109 33 121
rect 63 497 129 509
rect 63 121 79 497
rect 113 121 129 497
rect 63 109 129 121
rect 159 497 225 509
rect 159 121 175 497
rect 209 121 225 497
rect 159 109 225 121
rect 255 497 321 509
rect 255 121 271 497
rect 305 121 321 497
rect 255 109 321 121
rect 351 497 417 509
rect 351 121 367 497
rect 401 121 417 497
rect 351 109 417 121
rect 447 497 513 509
rect 447 121 463 497
rect 497 121 513 497
rect 447 109 513 121
rect 543 497 609 509
rect 543 121 559 497
rect 593 121 609 497
rect 543 109 609 121
rect 639 497 705 509
rect 639 121 655 497
rect 689 121 705 497
rect 639 109 705 121
rect 735 497 801 509
rect 735 121 751 497
rect 785 121 801 497
rect 735 109 801 121
rect 831 497 897 509
rect 831 121 847 497
rect 881 121 897 497
rect 831 109 897 121
rect 927 497 993 509
rect 927 121 943 497
rect 977 121 993 497
rect 927 109 993 121
rect 1023 497 1089 509
rect 1023 121 1039 497
rect 1073 121 1089 497
rect 1023 109 1089 121
rect 1119 497 1185 509
rect 1119 121 1135 497
rect 1169 121 1185 497
rect 1119 109 1185 121
rect 1215 497 1281 509
rect 1215 121 1231 497
rect 1265 121 1281 497
rect 1215 109 1281 121
rect 1311 497 1377 509
rect 1311 121 1327 497
rect 1361 121 1377 497
rect 1311 109 1377 121
rect 1407 497 1473 509
rect 1407 121 1423 497
rect 1457 121 1473 497
rect 1407 109 1473 121
rect 1503 497 1569 509
rect 1503 121 1519 497
rect 1553 121 1569 497
rect 1503 109 1569 121
rect 1599 497 1665 509
rect 1599 121 1615 497
rect 1649 121 1665 497
rect 1599 109 1665 121
rect 1695 497 1761 509
rect 1695 121 1711 497
rect 1745 121 1761 497
rect 1695 109 1761 121
rect 1791 497 1857 509
rect 1791 121 1807 497
rect 1841 121 1857 497
rect 1791 109 1857 121
rect 1887 497 1953 509
rect 1887 121 1903 497
rect 1937 121 1953 497
rect 1887 109 1953 121
rect 1983 497 2049 509
rect 1983 121 1999 497
rect 2033 121 2049 497
rect 1983 109 2049 121
rect 2079 497 2145 509
rect 2079 121 2095 497
rect 2129 121 2145 497
rect 2079 109 2145 121
rect 2175 497 2241 509
rect 2175 121 2191 497
rect 2225 121 2241 497
rect 2175 109 2241 121
rect 2271 497 2337 509
rect 2271 121 2287 497
rect 2321 121 2337 497
rect 2271 109 2337 121
rect 2367 497 2429 509
rect 2367 121 2383 497
rect 2417 121 2429 497
rect 2367 109 2429 121
rect -2429 -121 -2367 -109
rect -2429 -497 -2417 -121
rect -2383 -497 -2367 -121
rect -2429 -509 -2367 -497
rect -2337 -121 -2271 -109
rect -2337 -497 -2321 -121
rect -2287 -497 -2271 -121
rect -2337 -509 -2271 -497
rect -2241 -121 -2175 -109
rect -2241 -497 -2225 -121
rect -2191 -497 -2175 -121
rect -2241 -509 -2175 -497
rect -2145 -121 -2079 -109
rect -2145 -497 -2129 -121
rect -2095 -497 -2079 -121
rect -2145 -509 -2079 -497
rect -2049 -121 -1983 -109
rect -2049 -497 -2033 -121
rect -1999 -497 -1983 -121
rect -2049 -509 -1983 -497
rect -1953 -121 -1887 -109
rect -1953 -497 -1937 -121
rect -1903 -497 -1887 -121
rect -1953 -509 -1887 -497
rect -1857 -121 -1791 -109
rect -1857 -497 -1841 -121
rect -1807 -497 -1791 -121
rect -1857 -509 -1791 -497
rect -1761 -121 -1695 -109
rect -1761 -497 -1745 -121
rect -1711 -497 -1695 -121
rect -1761 -509 -1695 -497
rect -1665 -121 -1599 -109
rect -1665 -497 -1649 -121
rect -1615 -497 -1599 -121
rect -1665 -509 -1599 -497
rect -1569 -121 -1503 -109
rect -1569 -497 -1553 -121
rect -1519 -497 -1503 -121
rect -1569 -509 -1503 -497
rect -1473 -121 -1407 -109
rect -1473 -497 -1457 -121
rect -1423 -497 -1407 -121
rect -1473 -509 -1407 -497
rect -1377 -121 -1311 -109
rect -1377 -497 -1361 -121
rect -1327 -497 -1311 -121
rect -1377 -509 -1311 -497
rect -1281 -121 -1215 -109
rect -1281 -497 -1265 -121
rect -1231 -497 -1215 -121
rect -1281 -509 -1215 -497
rect -1185 -121 -1119 -109
rect -1185 -497 -1169 -121
rect -1135 -497 -1119 -121
rect -1185 -509 -1119 -497
rect -1089 -121 -1023 -109
rect -1089 -497 -1073 -121
rect -1039 -497 -1023 -121
rect -1089 -509 -1023 -497
rect -993 -121 -927 -109
rect -993 -497 -977 -121
rect -943 -497 -927 -121
rect -993 -509 -927 -497
rect -897 -121 -831 -109
rect -897 -497 -881 -121
rect -847 -497 -831 -121
rect -897 -509 -831 -497
rect -801 -121 -735 -109
rect -801 -497 -785 -121
rect -751 -497 -735 -121
rect -801 -509 -735 -497
rect -705 -121 -639 -109
rect -705 -497 -689 -121
rect -655 -497 -639 -121
rect -705 -509 -639 -497
rect -609 -121 -543 -109
rect -609 -497 -593 -121
rect -559 -497 -543 -121
rect -609 -509 -543 -497
rect -513 -121 -447 -109
rect -513 -497 -497 -121
rect -463 -497 -447 -121
rect -513 -509 -447 -497
rect -417 -121 -351 -109
rect -417 -497 -401 -121
rect -367 -497 -351 -121
rect -417 -509 -351 -497
rect -321 -121 -255 -109
rect -321 -497 -305 -121
rect -271 -497 -255 -121
rect -321 -509 -255 -497
rect -225 -121 -159 -109
rect -225 -497 -209 -121
rect -175 -497 -159 -121
rect -225 -509 -159 -497
rect -129 -121 -63 -109
rect -129 -497 -113 -121
rect -79 -497 -63 -121
rect -129 -509 -63 -497
rect -33 -121 33 -109
rect -33 -497 -17 -121
rect 17 -497 33 -121
rect -33 -509 33 -497
rect 63 -121 129 -109
rect 63 -497 79 -121
rect 113 -497 129 -121
rect 63 -509 129 -497
rect 159 -121 225 -109
rect 159 -497 175 -121
rect 209 -497 225 -121
rect 159 -509 225 -497
rect 255 -121 321 -109
rect 255 -497 271 -121
rect 305 -497 321 -121
rect 255 -509 321 -497
rect 351 -121 417 -109
rect 351 -497 367 -121
rect 401 -497 417 -121
rect 351 -509 417 -497
rect 447 -121 513 -109
rect 447 -497 463 -121
rect 497 -497 513 -121
rect 447 -509 513 -497
rect 543 -121 609 -109
rect 543 -497 559 -121
rect 593 -497 609 -121
rect 543 -509 609 -497
rect 639 -121 705 -109
rect 639 -497 655 -121
rect 689 -497 705 -121
rect 639 -509 705 -497
rect 735 -121 801 -109
rect 735 -497 751 -121
rect 785 -497 801 -121
rect 735 -509 801 -497
rect 831 -121 897 -109
rect 831 -497 847 -121
rect 881 -497 897 -121
rect 831 -509 897 -497
rect 927 -121 993 -109
rect 927 -497 943 -121
rect 977 -497 993 -121
rect 927 -509 993 -497
rect 1023 -121 1089 -109
rect 1023 -497 1039 -121
rect 1073 -497 1089 -121
rect 1023 -509 1089 -497
rect 1119 -121 1185 -109
rect 1119 -497 1135 -121
rect 1169 -497 1185 -121
rect 1119 -509 1185 -497
rect 1215 -121 1281 -109
rect 1215 -497 1231 -121
rect 1265 -497 1281 -121
rect 1215 -509 1281 -497
rect 1311 -121 1377 -109
rect 1311 -497 1327 -121
rect 1361 -497 1377 -121
rect 1311 -509 1377 -497
rect 1407 -121 1473 -109
rect 1407 -497 1423 -121
rect 1457 -497 1473 -121
rect 1407 -509 1473 -497
rect 1503 -121 1569 -109
rect 1503 -497 1519 -121
rect 1553 -497 1569 -121
rect 1503 -509 1569 -497
rect 1599 -121 1665 -109
rect 1599 -497 1615 -121
rect 1649 -497 1665 -121
rect 1599 -509 1665 -497
rect 1695 -121 1761 -109
rect 1695 -497 1711 -121
rect 1745 -497 1761 -121
rect 1695 -509 1761 -497
rect 1791 -121 1857 -109
rect 1791 -497 1807 -121
rect 1841 -497 1857 -121
rect 1791 -509 1857 -497
rect 1887 -121 1953 -109
rect 1887 -497 1903 -121
rect 1937 -497 1953 -121
rect 1887 -509 1953 -497
rect 1983 -121 2049 -109
rect 1983 -497 1999 -121
rect 2033 -497 2049 -121
rect 1983 -509 2049 -497
rect 2079 -121 2145 -109
rect 2079 -497 2095 -121
rect 2129 -497 2145 -121
rect 2079 -509 2145 -497
rect 2175 -121 2241 -109
rect 2175 -497 2191 -121
rect 2225 -497 2241 -121
rect 2175 -509 2241 -497
rect 2271 -121 2337 -109
rect 2271 -497 2287 -121
rect 2321 -497 2337 -121
rect 2271 -509 2337 -497
rect 2367 -121 2429 -109
rect 2367 -497 2383 -121
rect 2417 -497 2429 -121
rect 2367 -509 2429 -497
<< ndiffc >>
rect -2417 121 -2383 497
rect -2321 121 -2287 497
rect -2225 121 -2191 497
rect -2129 121 -2095 497
rect -2033 121 -1999 497
rect -1937 121 -1903 497
rect -1841 121 -1807 497
rect -1745 121 -1711 497
rect -1649 121 -1615 497
rect -1553 121 -1519 497
rect -1457 121 -1423 497
rect -1361 121 -1327 497
rect -1265 121 -1231 497
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect 1231 121 1265 497
rect 1327 121 1361 497
rect 1423 121 1457 497
rect 1519 121 1553 497
rect 1615 121 1649 497
rect 1711 121 1745 497
rect 1807 121 1841 497
rect 1903 121 1937 497
rect 1999 121 2033 497
rect 2095 121 2129 497
rect 2191 121 2225 497
rect 2287 121 2321 497
rect 2383 121 2417 497
rect -2417 -497 -2383 -121
rect -2321 -497 -2287 -121
rect -2225 -497 -2191 -121
rect -2129 -497 -2095 -121
rect -2033 -497 -1999 -121
rect -1937 -497 -1903 -121
rect -1841 -497 -1807 -121
rect -1745 -497 -1711 -121
rect -1649 -497 -1615 -121
rect -1553 -497 -1519 -121
rect -1457 -497 -1423 -121
rect -1361 -497 -1327 -121
rect -1265 -497 -1231 -121
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect 1231 -497 1265 -121
rect 1327 -497 1361 -121
rect 1423 -497 1457 -121
rect 1519 -497 1553 -121
rect 1615 -497 1649 -121
rect 1711 -497 1745 -121
rect 1807 -497 1841 -121
rect 1903 -497 1937 -121
rect 1999 -497 2033 -121
rect 2095 -497 2129 -121
rect 2191 -497 2225 -121
rect 2287 -497 2321 -121
rect 2383 -497 2417 -121
<< psubdiff >>
rect -2531 649 -2435 683
rect 2435 649 2531 683
rect -2531 587 -2497 649
rect 2497 587 2531 649
rect -2531 -649 -2497 -587
rect 2497 -649 2531 -587
rect -2531 -683 -2435 -649
rect 2435 -683 2531 -649
<< psubdiffcont >>
rect -2435 649 2435 683
rect -2531 -587 -2497 587
rect 2497 -587 2531 587
rect -2435 -683 2435 -649
<< poly >>
rect -2385 581 -2319 597
rect -2385 547 -2369 581
rect -2335 547 -2319 581
rect -2385 531 -2319 547
rect -2193 581 -2127 597
rect -2193 547 -2177 581
rect -2143 547 -2127 581
rect -2367 509 -2337 531
rect -2271 509 -2241 535
rect -2193 531 -2127 547
rect -2001 581 -1935 597
rect -2001 547 -1985 581
rect -1951 547 -1935 581
rect -2175 509 -2145 531
rect -2079 509 -2049 535
rect -2001 531 -1935 547
rect -1809 581 -1743 597
rect -1809 547 -1793 581
rect -1759 547 -1743 581
rect -1983 509 -1953 531
rect -1887 509 -1857 535
rect -1809 531 -1743 547
rect -1617 581 -1551 597
rect -1617 547 -1601 581
rect -1567 547 -1551 581
rect -1791 509 -1761 531
rect -1695 509 -1665 535
rect -1617 531 -1551 547
rect -1425 581 -1359 597
rect -1425 547 -1409 581
rect -1375 547 -1359 581
rect -1599 509 -1569 531
rect -1503 509 -1473 535
rect -1425 531 -1359 547
rect -1233 581 -1167 597
rect -1233 547 -1217 581
rect -1183 547 -1167 581
rect -1407 509 -1377 531
rect -1311 509 -1281 535
rect -1233 531 -1167 547
rect -1041 581 -975 597
rect -1041 547 -1025 581
rect -991 547 -975 581
rect -1215 509 -1185 531
rect -1119 509 -1089 535
rect -1041 531 -975 547
rect -849 581 -783 597
rect -849 547 -833 581
rect -799 547 -783 581
rect -1023 509 -993 531
rect -927 509 -897 535
rect -849 531 -783 547
rect -657 581 -591 597
rect -657 547 -641 581
rect -607 547 -591 581
rect -831 509 -801 531
rect -735 509 -705 535
rect -657 531 -591 547
rect -465 581 -399 597
rect -465 547 -449 581
rect -415 547 -399 581
rect -639 509 -609 531
rect -543 509 -513 535
rect -465 531 -399 547
rect -273 581 -207 597
rect -273 547 -257 581
rect -223 547 -207 581
rect -447 509 -417 531
rect -351 509 -321 535
rect -273 531 -207 547
rect -81 581 -15 597
rect -81 547 -65 581
rect -31 547 -15 581
rect -255 509 -225 531
rect -159 509 -129 535
rect -81 531 -15 547
rect 111 581 177 597
rect 111 547 127 581
rect 161 547 177 581
rect -63 509 -33 531
rect 33 509 63 535
rect 111 531 177 547
rect 303 581 369 597
rect 303 547 319 581
rect 353 547 369 581
rect 129 509 159 531
rect 225 509 255 535
rect 303 531 369 547
rect 495 581 561 597
rect 495 547 511 581
rect 545 547 561 581
rect 321 509 351 531
rect 417 509 447 535
rect 495 531 561 547
rect 687 581 753 597
rect 687 547 703 581
rect 737 547 753 581
rect 513 509 543 531
rect 609 509 639 535
rect 687 531 753 547
rect 879 581 945 597
rect 879 547 895 581
rect 929 547 945 581
rect 705 509 735 531
rect 801 509 831 535
rect 879 531 945 547
rect 1071 581 1137 597
rect 1071 547 1087 581
rect 1121 547 1137 581
rect 897 509 927 531
rect 993 509 1023 535
rect 1071 531 1137 547
rect 1263 581 1329 597
rect 1263 547 1279 581
rect 1313 547 1329 581
rect 1089 509 1119 531
rect 1185 509 1215 535
rect 1263 531 1329 547
rect 1455 581 1521 597
rect 1455 547 1471 581
rect 1505 547 1521 581
rect 1281 509 1311 531
rect 1377 509 1407 535
rect 1455 531 1521 547
rect 1647 581 1713 597
rect 1647 547 1663 581
rect 1697 547 1713 581
rect 1473 509 1503 531
rect 1569 509 1599 535
rect 1647 531 1713 547
rect 1839 581 1905 597
rect 1839 547 1855 581
rect 1889 547 1905 581
rect 1665 509 1695 531
rect 1761 509 1791 535
rect 1839 531 1905 547
rect 2031 581 2097 597
rect 2031 547 2047 581
rect 2081 547 2097 581
rect 1857 509 1887 531
rect 1953 509 1983 535
rect 2031 531 2097 547
rect 2223 581 2289 597
rect 2223 547 2239 581
rect 2273 547 2289 581
rect 2049 509 2079 531
rect 2145 509 2175 535
rect 2223 531 2289 547
rect 2241 509 2271 531
rect 2337 509 2367 535
rect -2367 83 -2337 109
rect -2271 87 -2241 109
rect -2289 71 -2223 87
rect -2175 83 -2145 109
rect -2079 87 -2049 109
rect -2289 37 -2273 71
rect -2239 37 -2223 71
rect -2289 21 -2223 37
rect -2097 71 -2031 87
rect -1983 83 -1953 109
rect -1887 87 -1857 109
rect -2097 37 -2081 71
rect -2047 37 -2031 71
rect -2097 21 -2031 37
rect -1905 71 -1839 87
rect -1791 83 -1761 109
rect -1695 87 -1665 109
rect -1905 37 -1889 71
rect -1855 37 -1839 71
rect -1905 21 -1839 37
rect -1713 71 -1647 87
rect -1599 83 -1569 109
rect -1503 87 -1473 109
rect -1713 37 -1697 71
rect -1663 37 -1647 71
rect -1713 21 -1647 37
rect -1521 71 -1455 87
rect -1407 83 -1377 109
rect -1311 87 -1281 109
rect -1521 37 -1505 71
rect -1471 37 -1455 71
rect -1521 21 -1455 37
rect -1329 71 -1263 87
rect -1215 83 -1185 109
rect -1119 87 -1089 109
rect -1329 37 -1313 71
rect -1279 37 -1263 71
rect -1329 21 -1263 37
rect -1137 71 -1071 87
rect -1023 83 -993 109
rect -927 87 -897 109
rect -1137 37 -1121 71
rect -1087 37 -1071 71
rect -1137 21 -1071 37
rect -945 71 -879 87
rect -831 83 -801 109
rect -735 87 -705 109
rect -945 37 -929 71
rect -895 37 -879 71
rect -945 21 -879 37
rect -753 71 -687 87
rect -639 83 -609 109
rect -543 87 -513 109
rect -753 37 -737 71
rect -703 37 -687 71
rect -753 21 -687 37
rect -561 71 -495 87
rect -447 83 -417 109
rect -351 87 -321 109
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 513 83 543 109
rect 609 87 639 109
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect 591 71 657 87
rect 705 83 735 109
rect 801 87 831 109
rect 591 37 607 71
rect 641 37 657 71
rect 591 21 657 37
rect 783 71 849 87
rect 897 83 927 109
rect 993 87 1023 109
rect 783 37 799 71
rect 833 37 849 71
rect 783 21 849 37
rect 975 71 1041 87
rect 1089 83 1119 109
rect 1185 87 1215 109
rect 975 37 991 71
rect 1025 37 1041 71
rect 975 21 1041 37
rect 1167 71 1233 87
rect 1281 83 1311 109
rect 1377 87 1407 109
rect 1167 37 1183 71
rect 1217 37 1233 71
rect 1167 21 1233 37
rect 1359 71 1425 87
rect 1473 83 1503 109
rect 1569 87 1599 109
rect 1359 37 1375 71
rect 1409 37 1425 71
rect 1359 21 1425 37
rect 1551 71 1617 87
rect 1665 83 1695 109
rect 1761 87 1791 109
rect 1551 37 1567 71
rect 1601 37 1617 71
rect 1551 21 1617 37
rect 1743 71 1809 87
rect 1857 83 1887 109
rect 1953 87 1983 109
rect 1743 37 1759 71
rect 1793 37 1809 71
rect 1743 21 1809 37
rect 1935 71 2001 87
rect 2049 83 2079 109
rect 2145 87 2175 109
rect 1935 37 1951 71
rect 1985 37 2001 71
rect 1935 21 2001 37
rect 2127 71 2193 87
rect 2241 83 2271 109
rect 2337 87 2367 109
rect 2127 37 2143 71
rect 2177 37 2193 71
rect 2127 21 2193 37
rect 2319 71 2385 87
rect 2319 37 2335 71
rect 2369 37 2385 71
rect 2319 21 2385 37
rect -2289 -37 -2223 -21
rect -2289 -71 -2273 -37
rect -2239 -71 -2223 -37
rect -2367 -109 -2337 -83
rect -2289 -87 -2223 -71
rect -2097 -37 -2031 -21
rect -2097 -71 -2081 -37
rect -2047 -71 -2031 -37
rect -2271 -109 -2241 -87
rect -2175 -109 -2145 -83
rect -2097 -87 -2031 -71
rect -1905 -37 -1839 -21
rect -1905 -71 -1889 -37
rect -1855 -71 -1839 -37
rect -2079 -109 -2049 -87
rect -1983 -109 -1953 -83
rect -1905 -87 -1839 -71
rect -1713 -37 -1647 -21
rect -1713 -71 -1697 -37
rect -1663 -71 -1647 -37
rect -1887 -109 -1857 -87
rect -1791 -109 -1761 -83
rect -1713 -87 -1647 -71
rect -1521 -37 -1455 -21
rect -1521 -71 -1505 -37
rect -1471 -71 -1455 -37
rect -1695 -109 -1665 -87
rect -1599 -109 -1569 -83
rect -1521 -87 -1455 -71
rect -1329 -37 -1263 -21
rect -1329 -71 -1313 -37
rect -1279 -71 -1263 -37
rect -1503 -109 -1473 -87
rect -1407 -109 -1377 -83
rect -1329 -87 -1263 -71
rect -1137 -37 -1071 -21
rect -1137 -71 -1121 -37
rect -1087 -71 -1071 -37
rect -1311 -109 -1281 -87
rect -1215 -109 -1185 -83
rect -1137 -87 -1071 -71
rect -945 -37 -879 -21
rect -945 -71 -929 -37
rect -895 -71 -879 -37
rect -1119 -109 -1089 -87
rect -1023 -109 -993 -83
rect -945 -87 -879 -71
rect -753 -37 -687 -21
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -927 -109 -897 -87
rect -831 -109 -801 -83
rect -753 -87 -687 -71
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -735 -109 -705 -87
rect -639 -109 -609 -83
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -543 -109 -513 -87
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 591 -37 657 -21
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 417 -109 447 -87
rect 513 -109 543 -83
rect 591 -87 657 -71
rect 783 -37 849 -21
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 609 -109 639 -87
rect 705 -109 735 -83
rect 783 -87 849 -71
rect 975 -37 1041 -21
rect 975 -71 991 -37
rect 1025 -71 1041 -37
rect 801 -109 831 -87
rect 897 -109 927 -83
rect 975 -87 1041 -71
rect 1167 -37 1233 -21
rect 1167 -71 1183 -37
rect 1217 -71 1233 -37
rect 993 -109 1023 -87
rect 1089 -109 1119 -83
rect 1167 -87 1233 -71
rect 1359 -37 1425 -21
rect 1359 -71 1375 -37
rect 1409 -71 1425 -37
rect 1185 -109 1215 -87
rect 1281 -109 1311 -83
rect 1359 -87 1425 -71
rect 1551 -37 1617 -21
rect 1551 -71 1567 -37
rect 1601 -71 1617 -37
rect 1377 -109 1407 -87
rect 1473 -109 1503 -83
rect 1551 -87 1617 -71
rect 1743 -37 1809 -21
rect 1743 -71 1759 -37
rect 1793 -71 1809 -37
rect 1569 -109 1599 -87
rect 1665 -109 1695 -83
rect 1743 -87 1809 -71
rect 1935 -37 2001 -21
rect 1935 -71 1951 -37
rect 1985 -71 2001 -37
rect 1761 -109 1791 -87
rect 1857 -109 1887 -83
rect 1935 -87 2001 -71
rect 2127 -37 2193 -21
rect 2127 -71 2143 -37
rect 2177 -71 2193 -37
rect 1953 -109 1983 -87
rect 2049 -109 2079 -83
rect 2127 -87 2193 -71
rect 2319 -37 2385 -21
rect 2319 -71 2335 -37
rect 2369 -71 2385 -37
rect 2145 -109 2175 -87
rect 2241 -109 2271 -83
rect 2319 -87 2385 -71
rect 2337 -109 2367 -87
rect -2367 -531 -2337 -509
rect -2385 -547 -2319 -531
rect -2271 -535 -2241 -509
rect -2175 -531 -2145 -509
rect -2385 -581 -2369 -547
rect -2335 -581 -2319 -547
rect -2385 -597 -2319 -581
rect -2193 -547 -2127 -531
rect -2079 -535 -2049 -509
rect -1983 -531 -1953 -509
rect -2193 -581 -2177 -547
rect -2143 -581 -2127 -547
rect -2193 -597 -2127 -581
rect -2001 -547 -1935 -531
rect -1887 -535 -1857 -509
rect -1791 -531 -1761 -509
rect -2001 -581 -1985 -547
rect -1951 -581 -1935 -547
rect -2001 -597 -1935 -581
rect -1809 -547 -1743 -531
rect -1695 -535 -1665 -509
rect -1599 -531 -1569 -509
rect -1809 -581 -1793 -547
rect -1759 -581 -1743 -547
rect -1809 -597 -1743 -581
rect -1617 -547 -1551 -531
rect -1503 -535 -1473 -509
rect -1407 -531 -1377 -509
rect -1617 -581 -1601 -547
rect -1567 -581 -1551 -547
rect -1617 -597 -1551 -581
rect -1425 -547 -1359 -531
rect -1311 -535 -1281 -509
rect -1215 -531 -1185 -509
rect -1425 -581 -1409 -547
rect -1375 -581 -1359 -547
rect -1425 -597 -1359 -581
rect -1233 -547 -1167 -531
rect -1119 -535 -1089 -509
rect -1023 -531 -993 -509
rect -1233 -581 -1217 -547
rect -1183 -581 -1167 -547
rect -1233 -597 -1167 -581
rect -1041 -547 -975 -531
rect -927 -535 -897 -509
rect -831 -531 -801 -509
rect -1041 -581 -1025 -547
rect -991 -581 -975 -547
rect -1041 -597 -975 -581
rect -849 -547 -783 -531
rect -735 -535 -705 -509
rect -639 -531 -609 -509
rect -849 -581 -833 -547
rect -799 -581 -783 -547
rect -849 -597 -783 -581
rect -657 -547 -591 -531
rect -543 -535 -513 -509
rect -447 -531 -417 -509
rect -657 -581 -641 -547
rect -607 -581 -591 -547
rect -657 -597 -591 -581
rect -465 -547 -399 -531
rect -351 -535 -321 -509
rect -255 -531 -225 -509
rect -465 -581 -449 -547
rect -415 -581 -399 -547
rect -465 -597 -399 -581
rect -273 -547 -207 -531
rect -159 -535 -129 -509
rect -63 -531 -33 -509
rect -273 -581 -257 -547
rect -223 -581 -207 -547
rect -273 -597 -207 -581
rect -81 -547 -15 -531
rect 33 -535 63 -509
rect 129 -531 159 -509
rect -81 -581 -65 -547
rect -31 -581 -15 -547
rect -81 -597 -15 -581
rect 111 -547 177 -531
rect 225 -535 255 -509
rect 321 -531 351 -509
rect 111 -581 127 -547
rect 161 -581 177 -547
rect 111 -597 177 -581
rect 303 -547 369 -531
rect 417 -535 447 -509
rect 513 -531 543 -509
rect 303 -581 319 -547
rect 353 -581 369 -547
rect 303 -597 369 -581
rect 495 -547 561 -531
rect 609 -535 639 -509
rect 705 -531 735 -509
rect 495 -581 511 -547
rect 545 -581 561 -547
rect 495 -597 561 -581
rect 687 -547 753 -531
rect 801 -535 831 -509
rect 897 -531 927 -509
rect 687 -581 703 -547
rect 737 -581 753 -547
rect 687 -597 753 -581
rect 879 -547 945 -531
rect 993 -535 1023 -509
rect 1089 -531 1119 -509
rect 879 -581 895 -547
rect 929 -581 945 -547
rect 879 -597 945 -581
rect 1071 -547 1137 -531
rect 1185 -535 1215 -509
rect 1281 -531 1311 -509
rect 1071 -581 1087 -547
rect 1121 -581 1137 -547
rect 1071 -597 1137 -581
rect 1263 -547 1329 -531
rect 1377 -535 1407 -509
rect 1473 -531 1503 -509
rect 1263 -581 1279 -547
rect 1313 -581 1329 -547
rect 1263 -597 1329 -581
rect 1455 -547 1521 -531
rect 1569 -535 1599 -509
rect 1665 -531 1695 -509
rect 1455 -581 1471 -547
rect 1505 -581 1521 -547
rect 1455 -597 1521 -581
rect 1647 -547 1713 -531
rect 1761 -535 1791 -509
rect 1857 -531 1887 -509
rect 1647 -581 1663 -547
rect 1697 -581 1713 -547
rect 1647 -597 1713 -581
rect 1839 -547 1905 -531
rect 1953 -535 1983 -509
rect 2049 -531 2079 -509
rect 1839 -581 1855 -547
rect 1889 -581 1905 -547
rect 1839 -597 1905 -581
rect 2031 -547 2097 -531
rect 2145 -535 2175 -509
rect 2241 -531 2271 -509
rect 2031 -581 2047 -547
rect 2081 -581 2097 -547
rect 2031 -597 2097 -581
rect 2223 -547 2289 -531
rect 2337 -535 2367 -509
rect 2223 -581 2239 -547
rect 2273 -581 2289 -547
rect 2223 -597 2289 -581
<< polycont >>
rect -2369 547 -2335 581
rect -2177 547 -2143 581
rect -1985 547 -1951 581
rect -1793 547 -1759 581
rect -1601 547 -1567 581
rect -1409 547 -1375 581
rect -1217 547 -1183 581
rect -1025 547 -991 581
rect -833 547 -799 581
rect -641 547 -607 581
rect -449 547 -415 581
rect -257 547 -223 581
rect -65 547 -31 581
rect 127 547 161 581
rect 319 547 353 581
rect 511 547 545 581
rect 703 547 737 581
rect 895 547 929 581
rect 1087 547 1121 581
rect 1279 547 1313 581
rect 1471 547 1505 581
rect 1663 547 1697 581
rect 1855 547 1889 581
rect 2047 547 2081 581
rect 2239 547 2273 581
rect -2273 37 -2239 71
rect -2081 37 -2047 71
rect -1889 37 -1855 71
rect -1697 37 -1663 71
rect -1505 37 -1471 71
rect -1313 37 -1279 71
rect -1121 37 -1087 71
rect -929 37 -895 71
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect 991 37 1025 71
rect 1183 37 1217 71
rect 1375 37 1409 71
rect 1567 37 1601 71
rect 1759 37 1793 71
rect 1951 37 1985 71
rect 2143 37 2177 71
rect 2335 37 2369 71
rect -2273 -71 -2239 -37
rect -2081 -71 -2047 -37
rect -1889 -71 -1855 -37
rect -1697 -71 -1663 -37
rect -1505 -71 -1471 -37
rect -1313 -71 -1279 -37
rect -1121 -71 -1087 -37
rect -929 -71 -895 -37
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect 991 -71 1025 -37
rect 1183 -71 1217 -37
rect 1375 -71 1409 -37
rect 1567 -71 1601 -37
rect 1759 -71 1793 -37
rect 1951 -71 1985 -37
rect 2143 -71 2177 -37
rect 2335 -71 2369 -37
rect -2369 -581 -2335 -547
rect -2177 -581 -2143 -547
rect -1985 -581 -1951 -547
rect -1793 -581 -1759 -547
rect -1601 -581 -1567 -547
rect -1409 -581 -1375 -547
rect -1217 -581 -1183 -547
rect -1025 -581 -991 -547
rect -833 -581 -799 -547
rect -641 -581 -607 -547
rect -449 -581 -415 -547
rect -257 -581 -223 -547
rect -65 -581 -31 -547
rect 127 -581 161 -547
rect 319 -581 353 -547
rect 511 -581 545 -547
rect 703 -581 737 -547
rect 895 -581 929 -547
rect 1087 -581 1121 -547
rect 1279 -581 1313 -547
rect 1471 -581 1505 -547
rect 1663 -581 1697 -547
rect 1855 -581 1889 -547
rect 2047 -581 2081 -547
rect 2239 -581 2273 -547
<< locali >>
rect -2531 649 -2435 683
rect 2435 649 2531 683
rect -2531 587 -2497 649
rect 2497 587 2531 649
rect -2385 547 -2369 581
rect -2335 547 -2319 581
rect -2193 547 -2177 581
rect -2143 547 -2127 581
rect -2001 547 -1985 581
rect -1951 547 -1935 581
rect -1809 547 -1793 581
rect -1759 547 -1743 581
rect -1617 547 -1601 581
rect -1567 547 -1551 581
rect -1425 547 -1409 581
rect -1375 547 -1359 581
rect -1233 547 -1217 581
rect -1183 547 -1167 581
rect -1041 547 -1025 581
rect -991 547 -975 581
rect -849 547 -833 581
rect -799 547 -783 581
rect -657 547 -641 581
rect -607 547 -591 581
rect -465 547 -449 581
rect -415 547 -399 581
rect -273 547 -257 581
rect -223 547 -207 581
rect -81 547 -65 581
rect -31 547 -15 581
rect 111 547 127 581
rect 161 547 177 581
rect 303 547 319 581
rect 353 547 369 581
rect 495 547 511 581
rect 545 547 561 581
rect 687 547 703 581
rect 737 547 753 581
rect 879 547 895 581
rect 929 547 945 581
rect 1071 547 1087 581
rect 1121 547 1137 581
rect 1263 547 1279 581
rect 1313 547 1329 581
rect 1455 547 1471 581
rect 1505 547 1521 581
rect 1647 547 1663 581
rect 1697 547 1713 581
rect 1839 547 1855 581
rect 1889 547 1905 581
rect 2031 547 2047 581
rect 2081 547 2097 581
rect 2223 547 2239 581
rect 2273 547 2289 581
rect -2417 497 -2383 513
rect -2417 105 -2383 121
rect -2321 497 -2287 513
rect -2321 105 -2287 121
rect -2225 497 -2191 513
rect -2225 105 -2191 121
rect -2129 497 -2095 513
rect -2129 105 -2095 121
rect -2033 497 -1999 513
rect -2033 105 -1999 121
rect -1937 497 -1903 513
rect -1937 105 -1903 121
rect -1841 497 -1807 513
rect -1841 105 -1807 121
rect -1745 497 -1711 513
rect -1745 105 -1711 121
rect -1649 497 -1615 513
rect -1649 105 -1615 121
rect -1553 497 -1519 513
rect -1553 105 -1519 121
rect -1457 497 -1423 513
rect -1457 105 -1423 121
rect -1361 497 -1327 513
rect -1361 105 -1327 121
rect -1265 497 -1231 513
rect -1265 105 -1231 121
rect -1169 497 -1135 513
rect -1169 105 -1135 121
rect -1073 497 -1039 513
rect -1073 105 -1039 121
rect -977 497 -943 513
rect -977 105 -943 121
rect -881 497 -847 513
rect -881 105 -847 121
rect -785 497 -751 513
rect -785 105 -751 121
rect -689 497 -655 513
rect -689 105 -655 121
rect -593 497 -559 513
rect -593 105 -559 121
rect -497 497 -463 513
rect -497 105 -463 121
rect -401 497 -367 513
rect -401 105 -367 121
rect -305 497 -271 513
rect -305 105 -271 121
rect -209 497 -175 513
rect -209 105 -175 121
rect -113 497 -79 513
rect -113 105 -79 121
rect -17 497 17 513
rect -17 105 17 121
rect 79 497 113 513
rect 79 105 113 121
rect 175 497 209 513
rect 175 105 209 121
rect 271 497 305 513
rect 271 105 305 121
rect 367 497 401 513
rect 367 105 401 121
rect 463 497 497 513
rect 463 105 497 121
rect 559 497 593 513
rect 559 105 593 121
rect 655 497 689 513
rect 655 105 689 121
rect 751 497 785 513
rect 751 105 785 121
rect 847 497 881 513
rect 847 105 881 121
rect 943 497 977 513
rect 943 105 977 121
rect 1039 497 1073 513
rect 1039 105 1073 121
rect 1135 497 1169 513
rect 1135 105 1169 121
rect 1231 497 1265 513
rect 1231 105 1265 121
rect 1327 497 1361 513
rect 1327 105 1361 121
rect 1423 497 1457 513
rect 1423 105 1457 121
rect 1519 497 1553 513
rect 1519 105 1553 121
rect 1615 497 1649 513
rect 1615 105 1649 121
rect 1711 497 1745 513
rect 1711 105 1745 121
rect 1807 497 1841 513
rect 1807 105 1841 121
rect 1903 497 1937 513
rect 1903 105 1937 121
rect 1999 497 2033 513
rect 1999 105 2033 121
rect 2095 497 2129 513
rect 2095 105 2129 121
rect 2191 497 2225 513
rect 2191 105 2225 121
rect 2287 497 2321 513
rect 2287 105 2321 121
rect 2383 497 2417 513
rect 2383 105 2417 121
rect -2289 37 -2273 71
rect -2239 37 -2223 71
rect -2097 37 -2081 71
rect -2047 37 -2031 71
rect -1905 37 -1889 71
rect -1855 37 -1839 71
rect -1713 37 -1697 71
rect -1663 37 -1647 71
rect -1521 37 -1505 71
rect -1471 37 -1455 71
rect -1329 37 -1313 71
rect -1279 37 -1263 71
rect -1137 37 -1121 71
rect -1087 37 -1071 71
rect -945 37 -929 71
rect -895 37 -879 71
rect -753 37 -737 71
rect -703 37 -687 71
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect 591 37 607 71
rect 641 37 657 71
rect 783 37 799 71
rect 833 37 849 71
rect 975 37 991 71
rect 1025 37 1041 71
rect 1167 37 1183 71
rect 1217 37 1233 71
rect 1359 37 1375 71
rect 1409 37 1425 71
rect 1551 37 1567 71
rect 1601 37 1617 71
rect 1743 37 1759 71
rect 1793 37 1809 71
rect 1935 37 1951 71
rect 1985 37 2001 71
rect 2127 37 2143 71
rect 2177 37 2193 71
rect 2319 37 2335 71
rect 2369 37 2385 71
rect -2289 -71 -2273 -37
rect -2239 -71 -2223 -37
rect -2097 -71 -2081 -37
rect -2047 -71 -2031 -37
rect -1905 -71 -1889 -37
rect -1855 -71 -1839 -37
rect -1713 -71 -1697 -37
rect -1663 -71 -1647 -37
rect -1521 -71 -1505 -37
rect -1471 -71 -1455 -37
rect -1329 -71 -1313 -37
rect -1279 -71 -1263 -37
rect -1137 -71 -1121 -37
rect -1087 -71 -1071 -37
rect -945 -71 -929 -37
rect -895 -71 -879 -37
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 975 -71 991 -37
rect 1025 -71 1041 -37
rect 1167 -71 1183 -37
rect 1217 -71 1233 -37
rect 1359 -71 1375 -37
rect 1409 -71 1425 -37
rect 1551 -71 1567 -37
rect 1601 -71 1617 -37
rect 1743 -71 1759 -37
rect 1793 -71 1809 -37
rect 1935 -71 1951 -37
rect 1985 -71 2001 -37
rect 2127 -71 2143 -37
rect 2177 -71 2193 -37
rect 2319 -71 2335 -37
rect 2369 -71 2385 -37
rect -2417 -121 -2383 -105
rect -2417 -513 -2383 -497
rect -2321 -121 -2287 -105
rect -2321 -513 -2287 -497
rect -2225 -121 -2191 -105
rect -2225 -513 -2191 -497
rect -2129 -121 -2095 -105
rect -2129 -513 -2095 -497
rect -2033 -121 -1999 -105
rect -2033 -513 -1999 -497
rect -1937 -121 -1903 -105
rect -1937 -513 -1903 -497
rect -1841 -121 -1807 -105
rect -1841 -513 -1807 -497
rect -1745 -121 -1711 -105
rect -1745 -513 -1711 -497
rect -1649 -121 -1615 -105
rect -1649 -513 -1615 -497
rect -1553 -121 -1519 -105
rect -1553 -513 -1519 -497
rect -1457 -121 -1423 -105
rect -1457 -513 -1423 -497
rect -1361 -121 -1327 -105
rect -1361 -513 -1327 -497
rect -1265 -121 -1231 -105
rect -1265 -513 -1231 -497
rect -1169 -121 -1135 -105
rect -1169 -513 -1135 -497
rect -1073 -121 -1039 -105
rect -1073 -513 -1039 -497
rect -977 -121 -943 -105
rect -977 -513 -943 -497
rect -881 -121 -847 -105
rect -881 -513 -847 -497
rect -785 -121 -751 -105
rect -785 -513 -751 -497
rect -689 -121 -655 -105
rect -689 -513 -655 -497
rect -593 -121 -559 -105
rect -593 -513 -559 -497
rect -497 -121 -463 -105
rect -497 -513 -463 -497
rect -401 -121 -367 -105
rect -401 -513 -367 -497
rect -305 -121 -271 -105
rect -305 -513 -271 -497
rect -209 -121 -175 -105
rect -209 -513 -175 -497
rect -113 -121 -79 -105
rect -113 -513 -79 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 79 -121 113 -105
rect 79 -513 113 -497
rect 175 -121 209 -105
rect 175 -513 209 -497
rect 271 -121 305 -105
rect 271 -513 305 -497
rect 367 -121 401 -105
rect 367 -513 401 -497
rect 463 -121 497 -105
rect 463 -513 497 -497
rect 559 -121 593 -105
rect 559 -513 593 -497
rect 655 -121 689 -105
rect 655 -513 689 -497
rect 751 -121 785 -105
rect 751 -513 785 -497
rect 847 -121 881 -105
rect 847 -513 881 -497
rect 943 -121 977 -105
rect 943 -513 977 -497
rect 1039 -121 1073 -105
rect 1039 -513 1073 -497
rect 1135 -121 1169 -105
rect 1135 -513 1169 -497
rect 1231 -121 1265 -105
rect 1231 -513 1265 -497
rect 1327 -121 1361 -105
rect 1327 -513 1361 -497
rect 1423 -121 1457 -105
rect 1423 -513 1457 -497
rect 1519 -121 1553 -105
rect 1519 -513 1553 -497
rect 1615 -121 1649 -105
rect 1615 -513 1649 -497
rect 1711 -121 1745 -105
rect 1711 -513 1745 -497
rect 1807 -121 1841 -105
rect 1807 -513 1841 -497
rect 1903 -121 1937 -105
rect 1903 -513 1937 -497
rect 1999 -121 2033 -105
rect 1999 -513 2033 -497
rect 2095 -121 2129 -105
rect 2095 -513 2129 -497
rect 2191 -121 2225 -105
rect 2191 -513 2225 -497
rect 2287 -121 2321 -105
rect 2287 -513 2321 -497
rect 2383 -121 2417 -105
rect 2383 -513 2417 -497
rect -2385 -581 -2369 -547
rect -2335 -581 -2319 -547
rect -2193 -581 -2177 -547
rect -2143 -581 -2127 -547
rect -2001 -581 -1985 -547
rect -1951 -581 -1935 -547
rect -1809 -581 -1793 -547
rect -1759 -581 -1743 -547
rect -1617 -581 -1601 -547
rect -1567 -581 -1551 -547
rect -1425 -581 -1409 -547
rect -1375 -581 -1359 -547
rect -1233 -581 -1217 -547
rect -1183 -581 -1167 -547
rect -1041 -581 -1025 -547
rect -991 -581 -975 -547
rect -849 -581 -833 -547
rect -799 -581 -783 -547
rect -657 -581 -641 -547
rect -607 -581 -591 -547
rect -465 -581 -449 -547
rect -415 -581 -399 -547
rect -273 -581 -257 -547
rect -223 -581 -207 -547
rect -81 -581 -65 -547
rect -31 -581 -15 -547
rect 111 -581 127 -547
rect 161 -581 177 -547
rect 303 -581 319 -547
rect 353 -581 369 -547
rect 495 -581 511 -547
rect 545 -581 561 -547
rect 687 -581 703 -547
rect 737 -581 753 -547
rect 879 -581 895 -547
rect 929 -581 945 -547
rect 1071 -581 1087 -547
rect 1121 -581 1137 -547
rect 1263 -581 1279 -547
rect 1313 -581 1329 -547
rect 1455 -581 1471 -547
rect 1505 -581 1521 -547
rect 1647 -581 1663 -547
rect 1697 -581 1713 -547
rect 1839 -581 1855 -547
rect 1889 -581 1905 -547
rect 2031 -581 2047 -547
rect 2081 -581 2097 -547
rect 2223 -581 2239 -547
rect 2273 -581 2289 -547
rect -2531 -649 -2497 -587
rect 2497 -649 2531 -587
rect -2531 -683 -2435 -649
rect 2435 -683 2531 -649
<< viali >>
rect -2369 547 -2335 581
rect -2177 547 -2143 581
rect -1985 547 -1951 581
rect -1793 547 -1759 581
rect -1601 547 -1567 581
rect -1409 547 -1375 581
rect -1217 547 -1183 581
rect -1025 547 -991 581
rect -833 547 -799 581
rect -641 547 -607 581
rect -449 547 -415 581
rect -257 547 -223 581
rect -65 547 -31 581
rect 127 547 161 581
rect 319 547 353 581
rect 511 547 545 581
rect 703 547 737 581
rect 895 547 929 581
rect 1087 547 1121 581
rect 1279 547 1313 581
rect 1471 547 1505 581
rect 1663 547 1697 581
rect 1855 547 1889 581
rect 2047 547 2081 581
rect 2239 547 2273 581
rect -2417 121 -2383 497
rect -2321 121 -2287 497
rect -2225 121 -2191 497
rect -2129 121 -2095 497
rect -2033 121 -1999 497
rect -1937 121 -1903 497
rect -1841 121 -1807 497
rect -1745 121 -1711 497
rect -1649 121 -1615 497
rect -1553 121 -1519 497
rect -1457 121 -1423 497
rect -1361 121 -1327 497
rect -1265 121 -1231 497
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect 1231 121 1265 497
rect 1327 121 1361 497
rect 1423 121 1457 497
rect 1519 121 1553 497
rect 1615 121 1649 497
rect 1711 121 1745 497
rect 1807 121 1841 497
rect 1903 121 1937 497
rect 1999 121 2033 497
rect 2095 121 2129 497
rect 2191 121 2225 497
rect 2287 121 2321 497
rect 2383 121 2417 497
rect -2273 37 -2239 71
rect -2081 37 -2047 71
rect -1889 37 -1855 71
rect -1697 37 -1663 71
rect -1505 37 -1471 71
rect -1313 37 -1279 71
rect -1121 37 -1087 71
rect -929 37 -895 71
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect 991 37 1025 71
rect 1183 37 1217 71
rect 1375 37 1409 71
rect 1567 37 1601 71
rect 1759 37 1793 71
rect 1951 37 1985 71
rect 2143 37 2177 71
rect 2335 37 2369 71
rect -2273 -71 -2239 -37
rect -2081 -71 -2047 -37
rect -1889 -71 -1855 -37
rect -1697 -71 -1663 -37
rect -1505 -71 -1471 -37
rect -1313 -71 -1279 -37
rect -1121 -71 -1087 -37
rect -929 -71 -895 -37
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect 991 -71 1025 -37
rect 1183 -71 1217 -37
rect 1375 -71 1409 -37
rect 1567 -71 1601 -37
rect 1759 -71 1793 -37
rect 1951 -71 1985 -37
rect 2143 -71 2177 -37
rect 2335 -71 2369 -37
rect -2417 -497 -2383 -121
rect -2321 -497 -2287 -121
rect -2225 -497 -2191 -121
rect -2129 -497 -2095 -121
rect -2033 -497 -1999 -121
rect -1937 -497 -1903 -121
rect -1841 -497 -1807 -121
rect -1745 -497 -1711 -121
rect -1649 -497 -1615 -121
rect -1553 -497 -1519 -121
rect -1457 -497 -1423 -121
rect -1361 -497 -1327 -121
rect -1265 -497 -1231 -121
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect 1231 -497 1265 -121
rect 1327 -497 1361 -121
rect 1423 -497 1457 -121
rect 1519 -497 1553 -121
rect 1615 -497 1649 -121
rect 1711 -497 1745 -121
rect 1807 -497 1841 -121
rect 1903 -497 1937 -121
rect 1999 -497 2033 -121
rect 2095 -497 2129 -121
rect 2191 -497 2225 -121
rect 2287 -497 2321 -121
rect 2383 -497 2417 -121
rect -2369 -581 -2335 -547
rect -2177 -581 -2143 -547
rect -1985 -581 -1951 -547
rect -1793 -581 -1759 -547
rect -1601 -581 -1567 -547
rect -1409 -581 -1375 -547
rect -1217 -581 -1183 -547
rect -1025 -581 -991 -547
rect -833 -581 -799 -547
rect -641 -581 -607 -547
rect -449 -581 -415 -547
rect -257 -581 -223 -547
rect -65 -581 -31 -547
rect 127 -581 161 -547
rect 319 -581 353 -547
rect 511 -581 545 -547
rect 703 -581 737 -547
rect 895 -581 929 -547
rect 1087 -581 1121 -547
rect 1279 -581 1313 -547
rect 1471 -581 1505 -547
rect 1663 -581 1697 -547
rect 1855 -581 1889 -547
rect 2047 -581 2081 -547
rect 2239 -581 2273 -547
<< metal1 >>
rect -2381 581 -2323 587
rect -2381 547 -2369 581
rect -2335 547 -2323 581
rect -2381 541 -2323 547
rect -2189 581 -2131 587
rect -2189 547 -2177 581
rect -2143 547 -2131 581
rect -2189 541 -2131 547
rect -1997 581 -1939 587
rect -1997 547 -1985 581
rect -1951 547 -1939 581
rect -1997 541 -1939 547
rect -1805 581 -1747 587
rect -1805 547 -1793 581
rect -1759 547 -1747 581
rect -1805 541 -1747 547
rect -1613 581 -1555 587
rect -1613 547 -1601 581
rect -1567 547 -1555 581
rect -1613 541 -1555 547
rect -1421 581 -1363 587
rect -1421 547 -1409 581
rect -1375 547 -1363 581
rect -1421 541 -1363 547
rect -1229 581 -1171 587
rect -1229 547 -1217 581
rect -1183 547 -1171 581
rect -1229 541 -1171 547
rect -1037 581 -979 587
rect -1037 547 -1025 581
rect -991 547 -979 581
rect -1037 541 -979 547
rect -845 581 -787 587
rect -845 547 -833 581
rect -799 547 -787 581
rect -845 541 -787 547
rect -653 581 -595 587
rect -653 547 -641 581
rect -607 547 -595 581
rect -653 541 -595 547
rect -461 581 -403 587
rect -461 547 -449 581
rect -415 547 -403 581
rect -461 541 -403 547
rect -269 581 -211 587
rect -269 547 -257 581
rect -223 547 -211 581
rect -269 541 -211 547
rect -77 581 -19 587
rect -77 547 -65 581
rect -31 547 -19 581
rect -77 541 -19 547
rect 115 581 173 587
rect 115 547 127 581
rect 161 547 173 581
rect 115 541 173 547
rect 307 581 365 587
rect 307 547 319 581
rect 353 547 365 581
rect 307 541 365 547
rect 499 581 557 587
rect 499 547 511 581
rect 545 547 557 581
rect 499 541 557 547
rect 691 581 749 587
rect 691 547 703 581
rect 737 547 749 581
rect 691 541 749 547
rect 883 581 941 587
rect 883 547 895 581
rect 929 547 941 581
rect 883 541 941 547
rect 1075 581 1133 587
rect 1075 547 1087 581
rect 1121 547 1133 581
rect 1075 541 1133 547
rect 1267 581 1325 587
rect 1267 547 1279 581
rect 1313 547 1325 581
rect 1267 541 1325 547
rect 1459 581 1517 587
rect 1459 547 1471 581
rect 1505 547 1517 581
rect 1459 541 1517 547
rect 1651 581 1709 587
rect 1651 547 1663 581
rect 1697 547 1709 581
rect 1651 541 1709 547
rect 1843 581 1901 587
rect 1843 547 1855 581
rect 1889 547 1901 581
rect 1843 541 1901 547
rect 2035 581 2093 587
rect 2035 547 2047 581
rect 2081 547 2093 581
rect 2035 541 2093 547
rect 2227 581 2285 587
rect 2227 547 2239 581
rect 2273 547 2285 581
rect 2227 541 2285 547
rect -2423 497 -2377 509
rect -2423 121 -2417 497
rect -2383 121 -2377 497
rect -2423 109 -2377 121
rect -2327 497 -2281 509
rect -2327 121 -2321 497
rect -2287 121 -2281 497
rect -2327 109 -2281 121
rect -2231 497 -2185 509
rect -2231 121 -2225 497
rect -2191 121 -2185 497
rect -2231 109 -2185 121
rect -2135 497 -2089 509
rect -2135 121 -2129 497
rect -2095 121 -2089 497
rect -2135 109 -2089 121
rect -2039 497 -1993 509
rect -2039 121 -2033 497
rect -1999 121 -1993 497
rect -2039 109 -1993 121
rect -1943 497 -1897 509
rect -1943 121 -1937 497
rect -1903 121 -1897 497
rect -1943 109 -1897 121
rect -1847 497 -1801 509
rect -1847 121 -1841 497
rect -1807 121 -1801 497
rect -1847 109 -1801 121
rect -1751 497 -1705 509
rect -1751 121 -1745 497
rect -1711 121 -1705 497
rect -1751 109 -1705 121
rect -1655 497 -1609 509
rect -1655 121 -1649 497
rect -1615 121 -1609 497
rect -1655 109 -1609 121
rect -1559 497 -1513 509
rect -1559 121 -1553 497
rect -1519 121 -1513 497
rect -1559 109 -1513 121
rect -1463 497 -1417 509
rect -1463 121 -1457 497
rect -1423 121 -1417 497
rect -1463 109 -1417 121
rect -1367 497 -1321 509
rect -1367 121 -1361 497
rect -1327 121 -1321 497
rect -1367 109 -1321 121
rect -1271 497 -1225 509
rect -1271 121 -1265 497
rect -1231 121 -1225 497
rect -1271 109 -1225 121
rect -1175 497 -1129 509
rect -1175 121 -1169 497
rect -1135 121 -1129 497
rect -1175 109 -1129 121
rect -1079 497 -1033 509
rect -1079 121 -1073 497
rect -1039 121 -1033 497
rect -1079 109 -1033 121
rect -983 497 -937 509
rect -983 121 -977 497
rect -943 121 -937 497
rect -983 109 -937 121
rect -887 497 -841 509
rect -887 121 -881 497
rect -847 121 -841 497
rect -887 109 -841 121
rect -791 497 -745 509
rect -791 121 -785 497
rect -751 121 -745 497
rect -791 109 -745 121
rect -695 497 -649 509
rect -695 121 -689 497
rect -655 121 -649 497
rect -695 109 -649 121
rect -599 497 -553 509
rect -599 121 -593 497
rect -559 121 -553 497
rect -599 109 -553 121
rect -503 497 -457 509
rect -503 121 -497 497
rect -463 121 -457 497
rect -503 109 -457 121
rect -407 497 -361 509
rect -407 121 -401 497
rect -367 121 -361 497
rect -407 109 -361 121
rect -311 497 -265 509
rect -311 121 -305 497
rect -271 121 -265 497
rect -311 109 -265 121
rect -215 497 -169 509
rect -215 121 -209 497
rect -175 121 -169 497
rect -215 109 -169 121
rect -119 497 -73 509
rect -119 121 -113 497
rect -79 121 -73 497
rect -119 109 -73 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 73 497 119 509
rect 73 121 79 497
rect 113 121 119 497
rect 73 109 119 121
rect 169 497 215 509
rect 169 121 175 497
rect 209 121 215 497
rect 169 109 215 121
rect 265 497 311 509
rect 265 121 271 497
rect 305 121 311 497
rect 265 109 311 121
rect 361 497 407 509
rect 361 121 367 497
rect 401 121 407 497
rect 361 109 407 121
rect 457 497 503 509
rect 457 121 463 497
rect 497 121 503 497
rect 457 109 503 121
rect 553 497 599 509
rect 553 121 559 497
rect 593 121 599 497
rect 553 109 599 121
rect 649 497 695 509
rect 649 121 655 497
rect 689 121 695 497
rect 649 109 695 121
rect 745 497 791 509
rect 745 121 751 497
rect 785 121 791 497
rect 745 109 791 121
rect 841 497 887 509
rect 841 121 847 497
rect 881 121 887 497
rect 841 109 887 121
rect 937 497 983 509
rect 937 121 943 497
rect 977 121 983 497
rect 937 109 983 121
rect 1033 497 1079 509
rect 1033 121 1039 497
rect 1073 121 1079 497
rect 1033 109 1079 121
rect 1129 497 1175 509
rect 1129 121 1135 497
rect 1169 121 1175 497
rect 1129 109 1175 121
rect 1225 497 1271 509
rect 1225 121 1231 497
rect 1265 121 1271 497
rect 1225 109 1271 121
rect 1321 497 1367 509
rect 1321 121 1327 497
rect 1361 121 1367 497
rect 1321 109 1367 121
rect 1417 497 1463 509
rect 1417 121 1423 497
rect 1457 121 1463 497
rect 1417 109 1463 121
rect 1513 497 1559 509
rect 1513 121 1519 497
rect 1553 121 1559 497
rect 1513 109 1559 121
rect 1609 497 1655 509
rect 1609 121 1615 497
rect 1649 121 1655 497
rect 1609 109 1655 121
rect 1705 497 1751 509
rect 1705 121 1711 497
rect 1745 121 1751 497
rect 1705 109 1751 121
rect 1801 497 1847 509
rect 1801 121 1807 497
rect 1841 121 1847 497
rect 1801 109 1847 121
rect 1897 497 1943 509
rect 1897 121 1903 497
rect 1937 121 1943 497
rect 1897 109 1943 121
rect 1993 497 2039 509
rect 1993 121 1999 497
rect 2033 121 2039 497
rect 1993 109 2039 121
rect 2089 497 2135 509
rect 2089 121 2095 497
rect 2129 121 2135 497
rect 2089 109 2135 121
rect 2185 497 2231 509
rect 2185 121 2191 497
rect 2225 121 2231 497
rect 2185 109 2231 121
rect 2281 497 2327 509
rect 2281 121 2287 497
rect 2321 121 2327 497
rect 2281 109 2327 121
rect 2377 497 2423 509
rect 2377 121 2383 497
rect 2417 121 2423 497
rect 2377 109 2423 121
rect -2285 71 -2227 77
rect -2285 37 -2273 71
rect -2239 37 -2227 71
rect -2285 31 -2227 37
rect -2093 71 -2035 77
rect -2093 37 -2081 71
rect -2047 37 -2035 71
rect -2093 31 -2035 37
rect -1901 71 -1843 77
rect -1901 37 -1889 71
rect -1855 37 -1843 71
rect -1901 31 -1843 37
rect -1709 71 -1651 77
rect -1709 37 -1697 71
rect -1663 37 -1651 71
rect -1709 31 -1651 37
rect -1517 71 -1459 77
rect -1517 37 -1505 71
rect -1471 37 -1459 71
rect -1517 31 -1459 37
rect -1325 71 -1267 77
rect -1325 37 -1313 71
rect -1279 37 -1267 71
rect -1325 31 -1267 37
rect -1133 71 -1075 77
rect -1133 37 -1121 71
rect -1087 37 -1075 71
rect -1133 31 -1075 37
rect -941 71 -883 77
rect -941 37 -929 71
rect -895 37 -883 71
rect -941 31 -883 37
rect -749 71 -691 77
rect -749 37 -737 71
rect -703 37 -691 71
rect -749 31 -691 37
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect 595 71 653 77
rect 595 37 607 71
rect 641 37 653 71
rect 595 31 653 37
rect 787 71 845 77
rect 787 37 799 71
rect 833 37 845 71
rect 787 31 845 37
rect 979 71 1037 77
rect 979 37 991 71
rect 1025 37 1037 71
rect 979 31 1037 37
rect 1171 71 1229 77
rect 1171 37 1183 71
rect 1217 37 1229 71
rect 1171 31 1229 37
rect 1363 71 1421 77
rect 1363 37 1375 71
rect 1409 37 1421 71
rect 1363 31 1421 37
rect 1555 71 1613 77
rect 1555 37 1567 71
rect 1601 37 1613 71
rect 1555 31 1613 37
rect 1747 71 1805 77
rect 1747 37 1759 71
rect 1793 37 1805 71
rect 1747 31 1805 37
rect 1939 71 1997 77
rect 1939 37 1951 71
rect 1985 37 1997 71
rect 1939 31 1997 37
rect 2131 71 2189 77
rect 2131 37 2143 71
rect 2177 37 2189 71
rect 2131 31 2189 37
rect 2323 71 2381 77
rect 2323 37 2335 71
rect 2369 37 2381 71
rect 2323 31 2381 37
rect -2285 -37 -2227 -31
rect -2285 -71 -2273 -37
rect -2239 -71 -2227 -37
rect -2285 -77 -2227 -71
rect -2093 -37 -2035 -31
rect -2093 -71 -2081 -37
rect -2047 -71 -2035 -37
rect -2093 -77 -2035 -71
rect -1901 -37 -1843 -31
rect -1901 -71 -1889 -37
rect -1855 -71 -1843 -37
rect -1901 -77 -1843 -71
rect -1709 -37 -1651 -31
rect -1709 -71 -1697 -37
rect -1663 -71 -1651 -37
rect -1709 -77 -1651 -71
rect -1517 -37 -1459 -31
rect -1517 -71 -1505 -37
rect -1471 -71 -1459 -37
rect -1517 -77 -1459 -71
rect -1325 -37 -1267 -31
rect -1325 -71 -1313 -37
rect -1279 -71 -1267 -37
rect -1325 -77 -1267 -71
rect -1133 -37 -1075 -31
rect -1133 -71 -1121 -37
rect -1087 -71 -1075 -37
rect -1133 -77 -1075 -71
rect -941 -37 -883 -31
rect -941 -71 -929 -37
rect -895 -71 -883 -37
rect -941 -77 -883 -71
rect -749 -37 -691 -31
rect -749 -71 -737 -37
rect -703 -71 -691 -37
rect -749 -77 -691 -71
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect 595 -37 653 -31
rect 595 -71 607 -37
rect 641 -71 653 -37
rect 595 -77 653 -71
rect 787 -37 845 -31
rect 787 -71 799 -37
rect 833 -71 845 -37
rect 787 -77 845 -71
rect 979 -37 1037 -31
rect 979 -71 991 -37
rect 1025 -71 1037 -37
rect 979 -77 1037 -71
rect 1171 -37 1229 -31
rect 1171 -71 1183 -37
rect 1217 -71 1229 -37
rect 1171 -77 1229 -71
rect 1363 -37 1421 -31
rect 1363 -71 1375 -37
rect 1409 -71 1421 -37
rect 1363 -77 1421 -71
rect 1555 -37 1613 -31
rect 1555 -71 1567 -37
rect 1601 -71 1613 -37
rect 1555 -77 1613 -71
rect 1747 -37 1805 -31
rect 1747 -71 1759 -37
rect 1793 -71 1805 -37
rect 1747 -77 1805 -71
rect 1939 -37 1997 -31
rect 1939 -71 1951 -37
rect 1985 -71 1997 -37
rect 1939 -77 1997 -71
rect 2131 -37 2189 -31
rect 2131 -71 2143 -37
rect 2177 -71 2189 -37
rect 2131 -77 2189 -71
rect 2323 -37 2381 -31
rect 2323 -71 2335 -37
rect 2369 -71 2381 -37
rect 2323 -77 2381 -71
rect -2423 -121 -2377 -109
rect -2423 -497 -2417 -121
rect -2383 -497 -2377 -121
rect -2423 -509 -2377 -497
rect -2327 -121 -2281 -109
rect -2327 -497 -2321 -121
rect -2287 -497 -2281 -121
rect -2327 -509 -2281 -497
rect -2231 -121 -2185 -109
rect -2231 -497 -2225 -121
rect -2191 -497 -2185 -121
rect -2231 -509 -2185 -497
rect -2135 -121 -2089 -109
rect -2135 -497 -2129 -121
rect -2095 -497 -2089 -121
rect -2135 -509 -2089 -497
rect -2039 -121 -1993 -109
rect -2039 -497 -2033 -121
rect -1999 -497 -1993 -121
rect -2039 -509 -1993 -497
rect -1943 -121 -1897 -109
rect -1943 -497 -1937 -121
rect -1903 -497 -1897 -121
rect -1943 -509 -1897 -497
rect -1847 -121 -1801 -109
rect -1847 -497 -1841 -121
rect -1807 -497 -1801 -121
rect -1847 -509 -1801 -497
rect -1751 -121 -1705 -109
rect -1751 -497 -1745 -121
rect -1711 -497 -1705 -121
rect -1751 -509 -1705 -497
rect -1655 -121 -1609 -109
rect -1655 -497 -1649 -121
rect -1615 -497 -1609 -121
rect -1655 -509 -1609 -497
rect -1559 -121 -1513 -109
rect -1559 -497 -1553 -121
rect -1519 -497 -1513 -121
rect -1559 -509 -1513 -497
rect -1463 -121 -1417 -109
rect -1463 -497 -1457 -121
rect -1423 -497 -1417 -121
rect -1463 -509 -1417 -497
rect -1367 -121 -1321 -109
rect -1367 -497 -1361 -121
rect -1327 -497 -1321 -121
rect -1367 -509 -1321 -497
rect -1271 -121 -1225 -109
rect -1271 -497 -1265 -121
rect -1231 -497 -1225 -121
rect -1271 -509 -1225 -497
rect -1175 -121 -1129 -109
rect -1175 -497 -1169 -121
rect -1135 -497 -1129 -121
rect -1175 -509 -1129 -497
rect -1079 -121 -1033 -109
rect -1079 -497 -1073 -121
rect -1039 -497 -1033 -121
rect -1079 -509 -1033 -497
rect -983 -121 -937 -109
rect -983 -497 -977 -121
rect -943 -497 -937 -121
rect -983 -509 -937 -497
rect -887 -121 -841 -109
rect -887 -497 -881 -121
rect -847 -497 -841 -121
rect -887 -509 -841 -497
rect -791 -121 -745 -109
rect -791 -497 -785 -121
rect -751 -497 -745 -121
rect -791 -509 -745 -497
rect -695 -121 -649 -109
rect -695 -497 -689 -121
rect -655 -497 -649 -121
rect -695 -509 -649 -497
rect -599 -121 -553 -109
rect -599 -497 -593 -121
rect -559 -497 -553 -121
rect -599 -509 -553 -497
rect -503 -121 -457 -109
rect -503 -497 -497 -121
rect -463 -497 -457 -121
rect -503 -509 -457 -497
rect -407 -121 -361 -109
rect -407 -497 -401 -121
rect -367 -497 -361 -121
rect -407 -509 -361 -497
rect -311 -121 -265 -109
rect -311 -497 -305 -121
rect -271 -497 -265 -121
rect -311 -509 -265 -497
rect -215 -121 -169 -109
rect -215 -497 -209 -121
rect -175 -497 -169 -121
rect -215 -509 -169 -497
rect -119 -121 -73 -109
rect -119 -497 -113 -121
rect -79 -497 -73 -121
rect -119 -509 -73 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 73 -121 119 -109
rect 73 -497 79 -121
rect 113 -497 119 -121
rect 73 -509 119 -497
rect 169 -121 215 -109
rect 169 -497 175 -121
rect 209 -497 215 -121
rect 169 -509 215 -497
rect 265 -121 311 -109
rect 265 -497 271 -121
rect 305 -497 311 -121
rect 265 -509 311 -497
rect 361 -121 407 -109
rect 361 -497 367 -121
rect 401 -497 407 -121
rect 361 -509 407 -497
rect 457 -121 503 -109
rect 457 -497 463 -121
rect 497 -497 503 -121
rect 457 -509 503 -497
rect 553 -121 599 -109
rect 553 -497 559 -121
rect 593 -497 599 -121
rect 553 -509 599 -497
rect 649 -121 695 -109
rect 649 -497 655 -121
rect 689 -497 695 -121
rect 649 -509 695 -497
rect 745 -121 791 -109
rect 745 -497 751 -121
rect 785 -497 791 -121
rect 745 -509 791 -497
rect 841 -121 887 -109
rect 841 -497 847 -121
rect 881 -497 887 -121
rect 841 -509 887 -497
rect 937 -121 983 -109
rect 937 -497 943 -121
rect 977 -497 983 -121
rect 937 -509 983 -497
rect 1033 -121 1079 -109
rect 1033 -497 1039 -121
rect 1073 -497 1079 -121
rect 1033 -509 1079 -497
rect 1129 -121 1175 -109
rect 1129 -497 1135 -121
rect 1169 -497 1175 -121
rect 1129 -509 1175 -497
rect 1225 -121 1271 -109
rect 1225 -497 1231 -121
rect 1265 -497 1271 -121
rect 1225 -509 1271 -497
rect 1321 -121 1367 -109
rect 1321 -497 1327 -121
rect 1361 -497 1367 -121
rect 1321 -509 1367 -497
rect 1417 -121 1463 -109
rect 1417 -497 1423 -121
rect 1457 -497 1463 -121
rect 1417 -509 1463 -497
rect 1513 -121 1559 -109
rect 1513 -497 1519 -121
rect 1553 -497 1559 -121
rect 1513 -509 1559 -497
rect 1609 -121 1655 -109
rect 1609 -497 1615 -121
rect 1649 -497 1655 -121
rect 1609 -509 1655 -497
rect 1705 -121 1751 -109
rect 1705 -497 1711 -121
rect 1745 -497 1751 -121
rect 1705 -509 1751 -497
rect 1801 -121 1847 -109
rect 1801 -497 1807 -121
rect 1841 -497 1847 -121
rect 1801 -509 1847 -497
rect 1897 -121 1943 -109
rect 1897 -497 1903 -121
rect 1937 -497 1943 -121
rect 1897 -509 1943 -497
rect 1993 -121 2039 -109
rect 1993 -497 1999 -121
rect 2033 -497 2039 -121
rect 1993 -509 2039 -497
rect 2089 -121 2135 -109
rect 2089 -497 2095 -121
rect 2129 -497 2135 -121
rect 2089 -509 2135 -497
rect 2185 -121 2231 -109
rect 2185 -497 2191 -121
rect 2225 -497 2231 -121
rect 2185 -509 2231 -497
rect 2281 -121 2327 -109
rect 2281 -497 2287 -121
rect 2321 -497 2327 -121
rect 2281 -509 2327 -497
rect 2377 -121 2423 -109
rect 2377 -497 2383 -121
rect 2417 -497 2423 -121
rect 2377 -509 2423 -497
rect -2381 -547 -2323 -541
rect -2381 -581 -2369 -547
rect -2335 -581 -2323 -547
rect -2381 -587 -2323 -581
rect -2189 -547 -2131 -541
rect -2189 -581 -2177 -547
rect -2143 -581 -2131 -547
rect -2189 -587 -2131 -581
rect -1997 -547 -1939 -541
rect -1997 -581 -1985 -547
rect -1951 -581 -1939 -547
rect -1997 -587 -1939 -581
rect -1805 -547 -1747 -541
rect -1805 -581 -1793 -547
rect -1759 -581 -1747 -547
rect -1805 -587 -1747 -581
rect -1613 -547 -1555 -541
rect -1613 -581 -1601 -547
rect -1567 -581 -1555 -547
rect -1613 -587 -1555 -581
rect -1421 -547 -1363 -541
rect -1421 -581 -1409 -547
rect -1375 -581 -1363 -547
rect -1421 -587 -1363 -581
rect -1229 -547 -1171 -541
rect -1229 -581 -1217 -547
rect -1183 -581 -1171 -547
rect -1229 -587 -1171 -581
rect -1037 -547 -979 -541
rect -1037 -581 -1025 -547
rect -991 -581 -979 -547
rect -1037 -587 -979 -581
rect -845 -547 -787 -541
rect -845 -581 -833 -547
rect -799 -581 -787 -547
rect -845 -587 -787 -581
rect -653 -547 -595 -541
rect -653 -581 -641 -547
rect -607 -581 -595 -547
rect -653 -587 -595 -581
rect -461 -547 -403 -541
rect -461 -581 -449 -547
rect -415 -581 -403 -547
rect -461 -587 -403 -581
rect -269 -547 -211 -541
rect -269 -581 -257 -547
rect -223 -581 -211 -547
rect -269 -587 -211 -581
rect -77 -547 -19 -541
rect -77 -581 -65 -547
rect -31 -581 -19 -547
rect -77 -587 -19 -581
rect 115 -547 173 -541
rect 115 -581 127 -547
rect 161 -581 173 -547
rect 115 -587 173 -581
rect 307 -547 365 -541
rect 307 -581 319 -547
rect 353 -581 365 -547
rect 307 -587 365 -581
rect 499 -547 557 -541
rect 499 -581 511 -547
rect 545 -581 557 -547
rect 499 -587 557 -581
rect 691 -547 749 -541
rect 691 -581 703 -547
rect 737 -581 749 -547
rect 691 -587 749 -581
rect 883 -547 941 -541
rect 883 -581 895 -547
rect 929 -581 941 -547
rect 883 -587 941 -581
rect 1075 -547 1133 -541
rect 1075 -581 1087 -547
rect 1121 -581 1133 -547
rect 1075 -587 1133 -581
rect 1267 -547 1325 -541
rect 1267 -581 1279 -547
rect 1313 -581 1325 -547
rect 1267 -587 1325 -581
rect 1459 -547 1517 -541
rect 1459 -581 1471 -547
rect 1505 -581 1517 -547
rect 1459 -587 1517 -581
rect 1651 -547 1709 -541
rect 1651 -581 1663 -547
rect 1697 -581 1709 -547
rect 1651 -587 1709 -581
rect 1843 -547 1901 -541
rect 1843 -581 1855 -547
rect 1889 -581 1901 -547
rect 1843 -587 1901 -581
rect 2035 -547 2093 -541
rect 2035 -581 2047 -547
rect 2081 -581 2093 -547
rect 2035 -587 2093 -581
rect 2227 -547 2285 -541
rect 2227 -581 2239 -547
rect 2273 -581 2285 -547
rect 2227 -587 2285 -581
<< properties >>
string FIXED_BBOX -2514 -666 2514 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 2 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
