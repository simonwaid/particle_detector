magic
tech sky130A
timestamp 1654768133
<< metal1 >>
rect 25 3340 50 3510
rect 440 3480 605 3510
rect 570 3365 595 3480
rect 330 3340 600 3365
rect 25 2200 50 2370
rect 455 2340 620 2370
rect 570 2200 595 2340
rect 25 1060 50 1230
rect 450 1200 595 1230
rect 570 1060 595 1200
rect 455 60 595 90
<< metal2 >>
rect 75 4495 200 4500
rect 75 4390 200 4395
rect 620 4495 745 4500
rect 620 4390 745 4395
rect 430 4250 1065 4325
rect 75 3355 200 3360
rect 75 3250 200 3255
rect 460 3135 520 3540
rect 620 3355 745 3360
rect 620 3250 745 3255
rect 1005 3130 1065 3535
rect 75 2215 200 2220
rect 75 2110 200 2115
rect 460 1985 520 2390
rect 620 2215 745 2220
rect 620 2110 745 2115
rect 1005 2030 1065 2435
rect 75 1075 200 1080
rect 75 970 200 975
rect 460 840 520 1245
rect 620 1075 745 1080
rect 620 970 745 975
rect 1005 870 1065 1275
<< via2 >>
rect 75 4395 200 4495
rect 620 4395 745 4495
rect 75 3255 200 3355
rect 620 3255 745 3355
rect 75 2115 200 2215
rect 620 2115 745 2215
rect 75 975 200 1075
rect 620 975 745 1075
<< metal3 >>
rect 70 4495 960 4570
rect 70 4395 75 4495
rect 200 4395 620 4495
rect 745 4395 960 4495
rect 70 4390 960 4395
rect 70 3355 205 4390
rect 70 3255 75 3355
rect 200 3255 205 3355
rect 70 2215 205 3255
rect 70 2115 75 2215
rect 200 2115 205 2215
rect 70 1075 205 2115
rect 70 975 75 1075
rect 200 975 205 1075
rect 70 970 205 975
rect 295 330 440 4050
rect 615 3355 750 4390
rect 615 3255 620 3355
rect 745 3255 750 3355
rect 615 2215 750 3255
rect 615 2115 620 2215
rect 745 2115 750 2215
rect 615 1075 750 2115
rect 615 975 620 1075
rect 745 975 750 1075
rect 615 970 750 975
rect 840 330 985 4050
rect 295 220 985 330
use bias_curm_p  bias_curm_p_0
timestamp 1654768133
transform 1 0 5 0 1 455
box -5 -455 550 695
use bias_curm_p  bias_curm_p_1
timestamp 1654768133
transform 1 0 550 0 1 455
box -5 -455 550 695
use bias_curm_p  bias_curm_p_2
timestamp 1654768133
transform 1 0 5 0 1 1595
box -5 -455 550 695
use bias_curm_p  bias_curm_p_3
timestamp 1654768133
transform 1 0 550 0 1 1595
box -5 -455 550 695
use bias_curm_p  bias_curm_p_4
timestamp 1654768133
transform 1 0 550 0 1 2735
box -5 -455 550 695
use bias_curm_p  bias_curm_p_5
timestamp 1654768133
transform 1 0 5 0 1 2735
box -5 -455 550 695
use bias_curm_p  bias_curm_p_6
timestamp 1654768133
transform 1 0 550 0 1 3875
box -5 -455 550 695
use bias_curm_p  bias_curm_p_7
timestamp 1654768133
transform 1 0 5 0 1 3875
box -5 -455 550 695
<< end >>
