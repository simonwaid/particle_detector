* SPICE3 file created from isource.ext - technology: sky130A

.subckt isource VP I_ref VN
X0 VP VM8D sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 VN VM3G VM3D VN sky130_fd_pr__nfet_01v8 ad=9.9185e+13p pd=7.231e+08u as=0p ps=0u w=4e+06u l=6e+06u
X2 VM3D VM3G VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X3 VM3D VM3G VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X4 VN VM3G VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X5 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.552e+13p ps=1.0376e+08u w=4e+06u l=150000u
X6 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X11 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X12 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X16 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X17 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X21 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X22 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X23 I_ref VM22D isource_out_0/m1_16760_11560# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X24 isource_out_0/m1_16760_11560# VM22D I_ref VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X25 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X26 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X27 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X28 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X29 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X30 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X31 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X32 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X33 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X34 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X35 isource_out_0/isource_cmirror_0/m1_250_820# VM8D VM22D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X36 isource_out_0/isource_cmirror_0/m1_250_820# VM8D VM22D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X37 VP VM8D isource_out_0/isource_cmirror_0/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=6.2785e+13p pd=4.649e+08u as=0p ps=0u w=4e+06u l=1e+06u
X38 VP VM8D isource_out_0/isource_cmirror_0/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X39 isource_out_0/isource_cmirror_0/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X40 VP VM8D isource_out_0/isource_cmirror_0/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X41 VP VM8D isource_out_0/isource_cmirror_0/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X42 isource_out_0/isource_cmirror_0/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X43 VP VM8D isource_out_0/isource_cmirror_0/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X44 VP VM8D isource_out_0/isource_cmirror_0/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X45 isource_out_0/isource_cmirror_0/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X46 isource_out_0/isource_cmirror_0/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X47 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X48 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X49 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X50 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X51 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X52 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X53 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X54 VM22D isource_out_0/m1_16760_11560# VM3D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X55 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X56 VM3D isource_out_0/m1_16760_11560# VM22D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X57 isource_out_0/m1_22920_9140# isource_out_0/m1_16760_11560# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X58 VN isource_out_0/m1_24520_11560# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X59 isource_out_0/m1_22920_9140# isource_out_0/m1_23460_11560# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X60 isource_out_0/m1_24000_9140# isource_out_0/m1_23460_11560# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X61 isource_out_0/m1_24000_9140# isource_out_0/m1_24520_11560# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X62 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.75622e+14p ps=1.58256e+09u w=4e+06u l=150000u
X63 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X64 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X65 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X66 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X67 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X68 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X69 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X70 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X71 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X72 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X73 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X74 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X75 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X76 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X77 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X78 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X79 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X80 VP VM14D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X81 VN VM14D VP VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X82 VP VN isource_startup_0/m1_330_800# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X83 VM8D isource_startup_0/m1_330_800# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X84 VN VN isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X85 isource_startup_0/m1_330_800# VN VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X86 isource_startup_0/m1_330_800# VN VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X87 VN VN isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X88 VN VN isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X89 isource_startup_0/m1_330_800# VN VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X90 isource_startup_0/m1_330_800# VN VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X91 isource_startup_0/m1_330_800# VN VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X92 VN VN isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X93 VN VN isource_startup_0/m1_330_800# VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X94 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X95 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X96 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X97 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X98 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X99 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X100 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X101 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X102 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X103 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X104 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X105 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X106 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X107 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X108 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X109 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X110 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X111 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X112 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X113 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X114 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X115 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X116 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X117 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X118 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X119 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X120 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X121 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X122 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X123 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X124 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X125 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X126 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X127 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X128 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X129 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X130 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X131 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X132 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X133 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X134 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X135 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X136 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X137 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X138 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X139 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X140 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X141 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X142 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X143 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X144 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X145 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X146 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X147 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X148 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X149 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X150 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X151 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X152 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X153 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X154 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X155 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X156 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X157 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X158 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X159 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X160 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X161 VN VM2D VM2D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X162 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X163 VM2D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X164 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X165 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X166 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X167 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X168 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X169 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X170 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X171 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X172 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X173 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X174 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X175 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X176 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X177 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X178 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X179 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X180 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X181 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X182 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X183 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X184 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X185 VM12D VM2D VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X186 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X187 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X188 VN VM2D VM12D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X189 VM12D VN isource_ref_0/sky130_fd_pr__nfet_01v8_WY4VMC_0/a_n1287_n400# isource_ref_0/sky130_fd_pr__nfet_01v8_WY4VMC_0/a_n1389_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X190 VN VN VM12D isource_ref_0/sky130_fd_pr__nfet_01v8_WY4VMC_0/a_n1389_n574# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X191 isource_cmirror_2/m1_250_820# VM8D VM9D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X192 isource_cmirror_2/m1_250_820# VM8D VM9D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X193 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X194 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X195 isource_cmirror_2/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X196 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X197 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X198 isource_cmirror_2/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X199 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X200 VP VM8D isource_cmirror_2/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X201 isource_cmirror_2/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X202 isource_cmirror_2/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X203 isource_cmirror_3/m1_250_820# VM8D VM8D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X204 isource_cmirror_3/m1_250_820# VM8D VM8D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X205 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X206 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X207 isource_cmirror_3/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X208 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X209 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X210 isource_cmirror_3/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X211 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X212 VP VM8D isource_cmirror_3/m1_250_820# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X213 isource_cmirror_3/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X214 isource_cmirror_3/m1_250_820# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X215 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X216 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X217 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X218 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X219 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X220 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X221 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X222 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X223 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X224 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X225 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X226 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X227 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X228 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X229 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X230 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X231 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X232 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X233 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X234 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X235 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X236 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X237 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X238 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X239 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X240 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X241 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X242 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X243 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X244 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X245 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X246 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X247 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X248 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X249 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X250 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X251 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X252 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X253 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X254 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X255 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X256 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X257 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X258 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X259 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X260 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X261 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X262 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X263 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X264 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X265 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X266 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X267 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X268 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X269 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X270 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X271 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X272 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X273 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X274 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X275 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X276 m2_19160_1520# VM8D VM14D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=200000u
X277 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X278 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X279 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X280 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X281 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X282 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X283 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X284 VP VM8D m2_19160_1520# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X285 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X286 m2_19160_1520# VM8D VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X287 isource_conv_0/m1_7960_7820# isource_conv_0/m1_7420_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X288 isource_conv_0/m1_6900_7820# isource_conv_0/m1_7420_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X289 VM3G isource_conv_0/m1_5300_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X290 isource_conv_0/m1_5840_7820# isource_conv_0/m1_5300_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X291 isource_conv_0/m1_5840_7820# isource_conv_0/m1_6360_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X292 VN isource_conv_0/m1_8480_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X293 isource_conv_0/m1_6900_7820# isource_conv_0/m1_6360_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X294 isource_conv_0/m1_7960_7820# isource_conv_0/m1_8480_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X295 VM14D VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X296 VN VN VM14D VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=6e+06u
X297 VM3G isource_conv_0/m1_4160_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X298 VN isource_conv_0/m1_4160_10260# VN sky130_fd_pr__res_xhigh_po_1p41 l=1e+07u
X299 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X300 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X301 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X302 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X303 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X304 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X305 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X306 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X307 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X308 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X309 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X310 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X311 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X312 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X313 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X314 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X315 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X316 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X317 VN VM9D VM8D VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X318 VM8D VM9D VN VN sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X319 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X320 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X321 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X322 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X323 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X324 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X325 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X326 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X327 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X328 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X329 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X330 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X331 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X332 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X333 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X334 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X335 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X336 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X337 VM2D VM9D VM9D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X338 VM9D VM9D VM2D VM2D sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X339 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X340 VN VP sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends
