magic
tech sky130B
magscale 1 2
timestamp 1654074216
<< pwell >>
rect -483 -719 483 719
<< nmos >>
rect -287 109 -187 509
rect -129 109 -29 509
rect 29 109 129 509
rect 187 109 287 509
rect -287 -509 -187 -109
rect -129 -509 -29 -109
rect 29 -509 129 -109
rect 187 -509 287 -109
<< ndiff >>
rect -345 497 -287 509
rect -345 121 -333 497
rect -299 121 -287 497
rect -345 109 -287 121
rect -187 497 -129 509
rect -187 121 -175 497
rect -141 121 -129 497
rect -187 109 -129 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 129 497 187 509
rect 129 121 141 497
rect 175 121 187 497
rect 129 109 187 121
rect 287 497 345 509
rect 287 121 299 497
rect 333 121 345 497
rect 287 109 345 121
rect -345 -121 -287 -109
rect -345 -497 -333 -121
rect -299 -497 -287 -121
rect -345 -509 -287 -497
rect -187 -121 -129 -109
rect -187 -497 -175 -121
rect -141 -497 -129 -121
rect -187 -509 -129 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 129 -121 187 -109
rect 129 -497 141 -121
rect 175 -497 187 -121
rect 129 -509 187 -497
rect 287 -121 345 -109
rect 287 -497 299 -121
rect 333 -497 345 -121
rect 287 -509 345 -497
<< ndiffc >>
rect -333 121 -299 497
rect -175 121 -141 497
rect -17 121 17 497
rect 141 121 175 497
rect 299 121 333 497
rect -333 -497 -299 -121
rect -175 -497 -141 -121
rect -17 -497 17 -121
rect 141 -497 175 -121
rect 299 -497 333 -121
<< psubdiff >>
rect -447 649 -351 683
rect 351 649 447 683
rect -447 587 -413 649
rect 413 587 447 649
rect -447 -649 -413 -587
rect 413 -649 447 -587
rect -447 -683 -351 -649
rect 351 -683 447 -649
<< psubdiffcont >>
rect -351 649 351 683
rect -447 -587 -413 587
rect 413 -587 447 587
rect -351 -683 351 -649
<< poly >>
rect -287 581 -187 597
rect -287 547 -271 581
rect -203 547 -187 581
rect -287 509 -187 547
rect -129 581 -29 597
rect -129 547 -113 581
rect -45 547 -29 581
rect -129 509 -29 547
rect 29 581 129 597
rect 29 547 45 581
rect 113 547 129 581
rect 29 509 129 547
rect 187 581 287 597
rect 187 547 203 581
rect 271 547 287 581
rect 187 509 287 547
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect -287 -547 -187 -509
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -287 -597 -187 -581
rect -129 -547 -29 -509
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -509
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 29 -597 129 -581
rect 187 -547 287 -509
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 187 -597 287 -581
<< polycont >>
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
<< locali >>
rect -447 649 -351 683
rect 351 649 447 683
rect -447 587 -413 649
rect 413 587 447 649
rect -287 547 -271 581
rect -203 547 -187 581
rect -129 547 -113 581
rect -45 547 -29 581
rect 29 547 45 581
rect 113 547 129 581
rect 187 547 203 581
rect 271 547 287 581
rect -333 497 -299 513
rect -333 105 -299 121
rect -175 497 -141 513
rect -175 105 -141 121
rect -17 497 17 513
rect -17 105 17 121
rect 141 497 175 513
rect 141 105 175 121
rect 299 497 333 513
rect 299 105 333 121
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect -333 -121 -299 -105
rect -333 -513 -299 -497
rect -175 -121 -141 -105
rect -175 -513 -141 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 141 -121 175 -105
rect 141 -513 175 -497
rect 299 -121 333 -105
rect 299 -513 333 -497
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 187 -581 203 -547
rect 271 -581 287 -547
rect -447 -649 -413 -587
rect 413 -649 447 -587
rect -447 -683 -351 -649
rect 351 -683 447 -649
<< viali >>
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect -333 121 -299 497
rect -175 121 -141 497
rect -17 121 17 497
rect 141 121 175 497
rect 299 121 333 497
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect -333 -497 -299 -121
rect -175 -497 -141 -121
rect -17 -497 17 -121
rect 141 -497 175 -121
rect 299 -497 333 -121
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
<< metal1 >>
rect -283 581 -191 587
rect -283 547 -271 581
rect -203 547 -191 581
rect -283 541 -191 547
rect -125 581 -33 587
rect -125 547 -113 581
rect -45 547 -33 581
rect -125 541 -33 547
rect 33 581 125 587
rect 33 547 45 581
rect 113 547 125 581
rect 33 541 125 547
rect 191 581 283 587
rect 191 547 203 581
rect 271 547 283 581
rect 191 541 283 547
rect -339 497 -293 509
rect -339 121 -333 497
rect -299 121 -293 497
rect -339 109 -293 121
rect -181 497 -135 509
rect -181 121 -175 497
rect -141 121 -135 497
rect -181 109 -135 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 135 497 181 509
rect 135 121 141 497
rect 175 121 181 497
rect 135 109 181 121
rect 293 497 339 509
rect 293 121 299 497
rect 333 121 339 497
rect 293 109 339 121
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect -339 -121 -293 -109
rect -339 -497 -333 -121
rect -299 -497 -293 -121
rect -339 -509 -293 -497
rect -181 -121 -135 -109
rect -181 -497 -175 -121
rect -141 -497 -135 -121
rect -181 -509 -135 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 135 -121 181 -109
rect 135 -497 141 -121
rect 175 -497 181 -121
rect 135 -509 181 -497
rect 293 -121 339 -109
rect 293 -497 299 -121
rect 333 -497 339 -121
rect 293 -509 339 -497
rect -283 -547 -191 -541
rect -283 -581 -271 -547
rect -203 -581 -191 -547
rect -283 -587 -191 -581
rect -125 -547 -33 -541
rect -125 -581 -113 -547
rect -45 -581 -33 -547
rect -125 -587 -33 -581
rect 33 -547 125 -541
rect 33 -581 45 -547
rect 113 -581 125 -547
rect 33 -587 125 -581
rect 191 -547 283 -541
rect 191 -581 203 -547
rect 271 -581 283 -547
rect 191 -587 283 -581
<< properties >>
string FIXED_BBOX -430 -666 430 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.5 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
