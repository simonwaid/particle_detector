magic
tech sky130A
magscale 1 2
timestamp 1645531774
<< nwell >>
rect -9073 127 -8407 1309
rect -8153 127 -7487 1309
rect -7233 127 -6567 1309
rect -6313 127 -5647 1309
rect -5393 127 -4727 1309
rect -4473 127 -3807 1309
rect -3553 127 -2887 1309
rect -2633 127 -1967 1309
rect -1713 127 -1047 1309
rect -793 127 -127 1309
rect 127 127 793 1309
rect 1047 127 1713 1309
rect 1967 127 2633 1309
rect 2887 127 3553 1309
rect 3807 127 4473 1309
rect 4727 127 5393 1309
rect 5647 127 6313 1309
rect 6567 127 7233 1309
rect 7487 127 8153 1309
rect 8407 127 9073 1309
rect -9073 -1309 -8407 -127
rect -8153 -1309 -7487 -127
rect -7233 -1309 -6567 -127
rect -6313 -1309 -5647 -127
rect -5393 -1309 -4727 -127
rect -4473 -1309 -3807 -127
rect -3553 -1309 -2887 -127
rect -2633 -1309 -1967 -127
rect -1713 -1309 -1047 -127
rect -793 -1309 -127 -127
rect 127 -1309 793 -127
rect 1047 -1309 1713 -127
rect 1967 -1309 2633 -127
rect 2887 -1309 3553 -127
rect 3807 -1309 4473 -127
rect 4727 -1309 5393 -127
rect 5647 -1309 6313 -127
rect 6567 -1309 7233 -127
rect 7487 -1309 8153 -127
rect 8407 -1309 9073 -127
<< pwell >>
rect -9183 1309 9183 1419
rect -9183 127 -9073 1309
rect -8407 127 -8153 1309
rect -7487 127 -7233 1309
rect -6567 127 -6313 1309
rect -5647 127 -5393 1309
rect -4727 127 -4473 1309
rect -3807 127 -3553 1309
rect -2887 127 -2633 1309
rect -1967 127 -1713 1309
rect -1047 127 -793 1309
rect -127 127 127 1309
rect 793 127 1047 1309
rect 1713 127 1967 1309
rect 2633 127 2887 1309
rect 3553 127 3807 1309
rect 4473 127 4727 1309
rect 5393 127 5647 1309
rect 6313 127 6567 1309
rect 7233 127 7487 1309
rect 8153 127 8407 1309
rect 9073 127 9183 1309
rect -9183 -127 9183 127
rect -9183 -1309 -9073 -127
rect -8407 -1309 -8153 -127
rect -7487 -1309 -7233 -127
rect -6567 -1309 -6313 -127
rect -5647 -1309 -5393 -127
rect -4727 -1309 -4473 -127
rect -3807 -1309 -3553 -127
rect -2887 -1309 -2633 -127
rect -1967 -1309 -1713 -127
rect -1047 -1309 -793 -127
rect -127 -1309 127 -127
rect 793 -1309 1047 -127
rect 1713 -1309 1967 -127
rect 2633 -1309 2887 -127
rect 3553 -1309 3807 -127
rect 4473 -1309 4727 -127
rect 5393 -1309 5647 -127
rect 6313 -1309 6567 -127
rect 7233 -1309 7487 -127
rect 8153 -1309 8407 -127
rect 9073 -1309 9183 -127
rect -9183 -1419 9183 -1309
<< varactor >>
rect -8940 218 -8540 1218
rect -8020 218 -7620 1218
rect -7100 218 -6700 1218
rect -6180 218 -5780 1218
rect -5260 218 -4860 1218
rect -4340 218 -3940 1218
rect -3420 218 -3020 1218
rect -2500 218 -2100 1218
rect -1580 218 -1180 1218
rect -660 218 -260 1218
rect 260 218 660 1218
rect 1180 218 1580 1218
rect 2100 218 2500 1218
rect 3020 218 3420 1218
rect 3940 218 4340 1218
rect 4860 218 5260 1218
rect 5780 218 6180 1218
rect 6700 218 7100 1218
rect 7620 218 8020 1218
rect 8540 218 8940 1218
rect -8940 -1218 -8540 -218
rect -8020 -1218 -7620 -218
rect -7100 -1218 -6700 -218
rect -6180 -1218 -5780 -218
rect -5260 -1218 -4860 -218
rect -4340 -1218 -3940 -218
rect -3420 -1218 -3020 -218
rect -2500 -1218 -2100 -218
rect -1580 -1218 -1180 -218
rect -660 -1218 -260 -218
rect 260 -1218 660 -218
rect 1180 -1218 1580 -218
rect 2100 -1218 2500 -218
rect 3020 -1218 3420 -218
rect 3940 -1218 4340 -218
rect 4860 -1218 5260 -218
rect 5780 -1218 6180 -218
rect 6700 -1218 7100 -218
rect 7620 -1218 8020 -218
rect 8540 -1218 8940 -218
<< psubdiff >>
rect -9147 1349 -9051 1383
rect 9051 1349 9147 1383
rect -9147 1287 -9113 1349
rect 9113 1287 9147 1349
rect -9147 -1349 -9113 -1287
rect 9113 -1349 9147 -1287
rect -9147 -1383 -9051 -1349
rect 9051 -1383 9147 -1349
<< nsubdiff >>
rect -9037 1194 -8940 1218
rect -9037 242 -9025 1194
rect -8991 242 -8940 1194
rect -9037 218 -8940 242
rect -8540 1194 -8443 1218
rect -8540 242 -8489 1194
rect -8455 242 -8443 1194
rect -8540 218 -8443 242
rect -8117 1194 -8020 1218
rect -8117 242 -8105 1194
rect -8071 242 -8020 1194
rect -8117 218 -8020 242
rect -7620 1194 -7523 1218
rect -7620 242 -7569 1194
rect -7535 242 -7523 1194
rect -7620 218 -7523 242
rect -7197 1194 -7100 1218
rect -7197 242 -7185 1194
rect -7151 242 -7100 1194
rect -7197 218 -7100 242
rect -6700 1194 -6603 1218
rect -6700 242 -6649 1194
rect -6615 242 -6603 1194
rect -6700 218 -6603 242
rect -6277 1194 -6180 1218
rect -6277 242 -6265 1194
rect -6231 242 -6180 1194
rect -6277 218 -6180 242
rect -5780 1194 -5683 1218
rect -5780 242 -5729 1194
rect -5695 242 -5683 1194
rect -5780 218 -5683 242
rect -5357 1194 -5260 1218
rect -5357 242 -5345 1194
rect -5311 242 -5260 1194
rect -5357 218 -5260 242
rect -4860 1194 -4763 1218
rect -4860 242 -4809 1194
rect -4775 242 -4763 1194
rect -4860 218 -4763 242
rect -4437 1194 -4340 1218
rect -4437 242 -4425 1194
rect -4391 242 -4340 1194
rect -4437 218 -4340 242
rect -3940 1194 -3843 1218
rect -3940 242 -3889 1194
rect -3855 242 -3843 1194
rect -3940 218 -3843 242
rect -3517 1194 -3420 1218
rect -3517 242 -3505 1194
rect -3471 242 -3420 1194
rect -3517 218 -3420 242
rect -3020 1194 -2923 1218
rect -3020 242 -2969 1194
rect -2935 242 -2923 1194
rect -3020 218 -2923 242
rect -2597 1194 -2500 1218
rect -2597 242 -2585 1194
rect -2551 242 -2500 1194
rect -2597 218 -2500 242
rect -2100 1194 -2003 1218
rect -2100 242 -2049 1194
rect -2015 242 -2003 1194
rect -2100 218 -2003 242
rect -1677 1194 -1580 1218
rect -1677 242 -1665 1194
rect -1631 242 -1580 1194
rect -1677 218 -1580 242
rect -1180 1194 -1083 1218
rect -1180 242 -1129 1194
rect -1095 242 -1083 1194
rect -1180 218 -1083 242
rect -757 1194 -660 1218
rect -757 242 -745 1194
rect -711 242 -660 1194
rect -757 218 -660 242
rect -260 1194 -163 1218
rect -260 242 -209 1194
rect -175 242 -163 1194
rect -260 218 -163 242
rect 163 1194 260 1218
rect 163 242 175 1194
rect 209 242 260 1194
rect 163 218 260 242
rect 660 1194 757 1218
rect 660 242 711 1194
rect 745 242 757 1194
rect 660 218 757 242
rect 1083 1194 1180 1218
rect 1083 242 1095 1194
rect 1129 242 1180 1194
rect 1083 218 1180 242
rect 1580 1194 1677 1218
rect 1580 242 1631 1194
rect 1665 242 1677 1194
rect 1580 218 1677 242
rect 2003 1194 2100 1218
rect 2003 242 2015 1194
rect 2049 242 2100 1194
rect 2003 218 2100 242
rect 2500 1194 2597 1218
rect 2500 242 2551 1194
rect 2585 242 2597 1194
rect 2500 218 2597 242
rect 2923 1194 3020 1218
rect 2923 242 2935 1194
rect 2969 242 3020 1194
rect 2923 218 3020 242
rect 3420 1194 3517 1218
rect 3420 242 3471 1194
rect 3505 242 3517 1194
rect 3420 218 3517 242
rect 3843 1194 3940 1218
rect 3843 242 3855 1194
rect 3889 242 3940 1194
rect 3843 218 3940 242
rect 4340 1194 4437 1218
rect 4340 242 4391 1194
rect 4425 242 4437 1194
rect 4340 218 4437 242
rect 4763 1194 4860 1218
rect 4763 242 4775 1194
rect 4809 242 4860 1194
rect 4763 218 4860 242
rect 5260 1194 5357 1218
rect 5260 242 5311 1194
rect 5345 242 5357 1194
rect 5260 218 5357 242
rect 5683 1194 5780 1218
rect 5683 242 5695 1194
rect 5729 242 5780 1194
rect 5683 218 5780 242
rect 6180 1194 6277 1218
rect 6180 242 6231 1194
rect 6265 242 6277 1194
rect 6180 218 6277 242
rect 6603 1194 6700 1218
rect 6603 242 6615 1194
rect 6649 242 6700 1194
rect 6603 218 6700 242
rect 7100 1194 7197 1218
rect 7100 242 7151 1194
rect 7185 242 7197 1194
rect 7100 218 7197 242
rect 7523 1194 7620 1218
rect 7523 242 7535 1194
rect 7569 242 7620 1194
rect 7523 218 7620 242
rect 8020 1194 8117 1218
rect 8020 242 8071 1194
rect 8105 242 8117 1194
rect 8020 218 8117 242
rect 8443 1194 8540 1218
rect 8443 242 8455 1194
rect 8489 242 8540 1194
rect 8443 218 8540 242
rect 8940 1194 9037 1218
rect 8940 242 8991 1194
rect 9025 242 9037 1194
rect 8940 218 9037 242
rect -9037 -242 -8940 -218
rect -9037 -1194 -9025 -242
rect -8991 -1194 -8940 -242
rect -9037 -1218 -8940 -1194
rect -8540 -242 -8443 -218
rect -8540 -1194 -8489 -242
rect -8455 -1194 -8443 -242
rect -8540 -1218 -8443 -1194
rect -8117 -242 -8020 -218
rect -8117 -1194 -8105 -242
rect -8071 -1194 -8020 -242
rect -8117 -1218 -8020 -1194
rect -7620 -242 -7523 -218
rect -7620 -1194 -7569 -242
rect -7535 -1194 -7523 -242
rect -7620 -1218 -7523 -1194
rect -7197 -242 -7100 -218
rect -7197 -1194 -7185 -242
rect -7151 -1194 -7100 -242
rect -7197 -1218 -7100 -1194
rect -6700 -242 -6603 -218
rect -6700 -1194 -6649 -242
rect -6615 -1194 -6603 -242
rect -6700 -1218 -6603 -1194
rect -6277 -242 -6180 -218
rect -6277 -1194 -6265 -242
rect -6231 -1194 -6180 -242
rect -6277 -1218 -6180 -1194
rect -5780 -242 -5683 -218
rect -5780 -1194 -5729 -242
rect -5695 -1194 -5683 -242
rect -5780 -1218 -5683 -1194
rect -5357 -242 -5260 -218
rect -5357 -1194 -5345 -242
rect -5311 -1194 -5260 -242
rect -5357 -1218 -5260 -1194
rect -4860 -242 -4763 -218
rect -4860 -1194 -4809 -242
rect -4775 -1194 -4763 -242
rect -4860 -1218 -4763 -1194
rect -4437 -242 -4340 -218
rect -4437 -1194 -4425 -242
rect -4391 -1194 -4340 -242
rect -4437 -1218 -4340 -1194
rect -3940 -242 -3843 -218
rect -3940 -1194 -3889 -242
rect -3855 -1194 -3843 -242
rect -3940 -1218 -3843 -1194
rect -3517 -242 -3420 -218
rect -3517 -1194 -3505 -242
rect -3471 -1194 -3420 -242
rect -3517 -1218 -3420 -1194
rect -3020 -242 -2923 -218
rect -3020 -1194 -2969 -242
rect -2935 -1194 -2923 -242
rect -3020 -1218 -2923 -1194
rect -2597 -242 -2500 -218
rect -2597 -1194 -2585 -242
rect -2551 -1194 -2500 -242
rect -2597 -1218 -2500 -1194
rect -2100 -242 -2003 -218
rect -2100 -1194 -2049 -242
rect -2015 -1194 -2003 -242
rect -2100 -1218 -2003 -1194
rect -1677 -242 -1580 -218
rect -1677 -1194 -1665 -242
rect -1631 -1194 -1580 -242
rect -1677 -1218 -1580 -1194
rect -1180 -242 -1083 -218
rect -1180 -1194 -1129 -242
rect -1095 -1194 -1083 -242
rect -1180 -1218 -1083 -1194
rect -757 -242 -660 -218
rect -757 -1194 -745 -242
rect -711 -1194 -660 -242
rect -757 -1218 -660 -1194
rect -260 -242 -163 -218
rect -260 -1194 -209 -242
rect -175 -1194 -163 -242
rect -260 -1218 -163 -1194
rect 163 -242 260 -218
rect 163 -1194 175 -242
rect 209 -1194 260 -242
rect 163 -1218 260 -1194
rect 660 -242 757 -218
rect 660 -1194 711 -242
rect 745 -1194 757 -242
rect 660 -1218 757 -1194
rect 1083 -242 1180 -218
rect 1083 -1194 1095 -242
rect 1129 -1194 1180 -242
rect 1083 -1218 1180 -1194
rect 1580 -242 1677 -218
rect 1580 -1194 1631 -242
rect 1665 -1194 1677 -242
rect 1580 -1218 1677 -1194
rect 2003 -242 2100 -218
rect 2003 -1194 2015 -242
rect 2049 -1194 2100 -242
rect 2003 -1218 2100 -1194
rect 2500 -242 2597 -218
rect 2500 -1194 2551 -242
rect 2585 -1194 2597 -242
rect 2500 -1218 2597 -1194
rect 2923 -242 3020 -218
rect 2923 -1194 2935 -242
rect 2969 -1194 3020 -242
rect 2923 -1218 3020 -1194
rect 3420 -242 3517 -218
rect 3420 -1194 3471 -242
rect 3505 -1194 3517 -242
rect 3420 -1218 3517 -1194
rect 3843 -242 3940 -218
rect 3843 -1194 3855 -242
rect 3889 -1194 3940 -242
rect 3843 -1218 3940 -1194
rect 4340 -242 4437 -218
rect 4340 -1194 4391 -242
rect 4425 -1194 4437 -242
rect 4340 -1218 4437 -1194
rect 4763 -242 4860 -218
rect 4763 -1194 4775 -242
rect 4809 -1194 4860 -242
rect 4763 -1218 4860 -1194
rect 5260 -242 5357 -218
rect 5260 -1194 5311 -242
rect 5345 -1194 5357 -242
rect 5260 -1218 5357 -1194
rect 5683 -242 5780 -218
rect 5683 -1194 5695 -242
rect 5729 -1194 5780 -242
rect 5683 -1218 5780 -1194
rect 6180 -242 6277 -218
rect 6180 -1194 6231 -242
rect 6265 -1194 6277 -242
rect 6180 -1218 6277 -1194
rect 6603 -242 6700 -218
rect 6603 -1194 6615 -242
rect 6649 -1194 6700 -242
rect 6603 -1218 6700 -1194
rect 7100 -242 7197 -218
rect 7100 -1194 7151 -242
rect 7185 -1194 7197 -242
rect 7100 -1218 7197 -1194
rect 7523 -242 7620 -218
rect 7523 -1194 7535 -242
rect 7569 -1194 7620 -242
rect 7523 -1218 7620 -1194
rect 8020 -242 8117 -218
rect 8020 -1194 8071 -242
rect 8105 -1194 8117 -242
rect 8020 -1218 8117 -1194
rect 8443 -242 8540 -218
rect 8443 -1194 8455 -242
rect 8489 -1194 8540 -242
rect 8443 -1218 8540 -1194
rect 8940 -242 9037 -218
rect 8940 -1194 8991 -242
rect 9025 -1194 9037 -242
rect 8940 -1218 9037 -1194
<< psubdiffcont >>
rect -9051 1349 9051 1383
rect -9147 -1287 -9113 1287
rect 9113 -1287 9147 1287
rect -9051 -1383 9051 -1349
<< nsubdiffcont >>
rect -9025 242 -8991 1194
rect -8489 242 -8455 1194
rect -8105 242 -8071 1194
rect -7569 242 -7535 1194
rect -7185 242 -7151 1194
rect -6649 242 -6615 1194
rect -6265 242 -6231 1194
rect -5729 242 -5695 1194
rect -5345 242 -5311 1194
rect -4809 242 -4775 1194
rect -4425 242 -4391 1194
rect -3889 242 -3855 1194
rect -3505 242 -3471 1194
rect -2969 242 -2935 1194
rect -2585 242 -2551 1194
rect -2049 242 -2015 1194
rect -1665 242 -1631 1194
rect -1129 242 -1095 1194
rect -745 242 -711 1194
rect -209 242 -175 1194
rect 175 242 209 1194
rect 711 242 745 1194
rect 1095 242 1129 1194
rect 1631 242 1665 1194
rect 2015 242 2049 1194
rect 2551 242 2585 1194
rect 2935 242 2969 1194
rect 3471 242 3505 1194
rect 3855 242 3889 1194
rect 4391 242 4425 1194
rect 4775 242 4809 1194
rect 5311 242 5345 1194
rect 5695 242 5729 1194
rect 6231 242 6265 1194
rect 6615 242 6649 1194
rect 7151 242 7185 1194
rect 7535 242 7569 1194
rect 8071 242 8105 1194
rect 8455 242 8489 1194
rect 8991 242 9025 1194
rect -9025 -1194 -8991 -242
rect -8489 -1194 -8455 -242
rect -8105 -1194 -8071 -242
rect -7569 -1194 -7535 -242
rect -7185 -1194 -7151 -242
rect -6649 -1194 -6615 -242
rect -6265 -1194 -6231 -242
rect -5729 -1194 -5695 -242
rect -5345 -1194 -5311 -242
rect -4809 -1194 -4775 -242
rect -4425 -1194 -4391 -242
rect -3889 -1194 -3855 -242
rect -3505 -1194 -3471 -242
rect -2969 -1194 -2935 -242
rect -2585 -1194 -2551 -242
rect -2049 -1194 -2015 -242
rect -1665 -1194 -1631 -242
rect -1129 -1194 -1095 -242
rect -745 -1194 -711 -242
rect -209 -1194 -175 -242
rect 175 -1194 209 -242
rect 711 -1194 745 -242
rect 1095 -1194 1129 -242
rect 1631 -1194 1665 -242
rect 2015 -1194 2049 -242
rect 2551 -1194 2585 -242
rect 2935 -1194 2969 -242
rect 3471 -1194 3505 -242
rect 3855 -1194 3889 -242
rect 4391 -1194 4425 -242
rect 4775 -1194 4809 -242
rect 5311 -1194 5345 -242
rect 5695 -1194 5729 -242
rect 6231 -1194 6265 -242
rect 6615 -1194 6649 -242
rect 7151 -1194 7185 -242
rect 7535 -1194 7569 -242
rect 8071 -1194 8105 -242
rect 8455 -1194 8489 -242
rect 8991 -1194 9025 -242
<< poly >>
rect -8940 1290 -8540 1306
rect -8940 1256 -8924 1290
rect -8556 1256 -8540 1290
rect -8940 1218 -8540 1256
rect -8020 1290 -7620 1306
rect -8020 1256 -8004 1290
rect -7636 1256 -7620 1290
rect -8020 1218 -7620 1256
rect -7100 1290 -6700 1306
rect -7100 1256 -7084 1290
rect -6716 1256 -6700 1290
rect -7100 1218 -6700 1256
rect -6180 1290 -5780 1306
rect -6180 1256 -6164 1290
rect -5796 1256 -5780 1290
rect -6180 1218 -5780 1256
rect -5260 1290 -4860 1306
rect -5260 1256 -5244 1290
rect -4876 1256 -4860 1290
rect -5260 1218 -4860 1256
rect -4340 1290 -3940 1306
rect -4340 1256 -4324 1290
rect -3956 1256 -3940 1290
rect -4340 1218 -3940 1256
rect -3420 1290 -3020 1306
rect -3420 1256 -3404 1290
rect -3036 1256 -3020 1290
rect -3420 1218 -3020 1256
rect -2500 1290 -2100 1306
rect -2500 1256 -2484 1290
rect -2116 1256 -2100 1290
rect -2500 1218 -2100 1256
rect -1580 1290 -1180 1306
rect -1580 1256 -1564 1290
rect -1196 1256 -1180 1290
rect -1580 1218 -1180 1256
rect -660 1290 -260 1306
rect -660 1256 -644 1290
rect -276 1256 -260 1290
rect -660 1218 -260 1256
rect 260 1290 660 1306
rect 260 1256 276 1290
rect 644 1256 660 1290
rect 260 1218 660 1256
rect 1180 1290 1580 1306
rect 1180 1256 1196 1290
rect 1564 1256 1580 1290
rect 1180 1218 1580 1256
rect 2100 1290 2500 1306
rect 2100 1256 2116 1290
rect 2484 1256 2500 1290
rect 2100 1218 2500 1256
rect 3020 1290 3420 1306
rect 3020 1256 3036 1290
rect 3404 1256 3420 1290
rect 3020 1218 3420 1256
rect 3940 1290 4340 1306
rect 3940 1256 3956 1290
rect 4324 1256 4340 1290
rect 3940 1218 4340 1256
rect 4860 1290 5260 1306
rect 4860 1256 4876 1290
rect 5244 1256 5260 1290
rect 4860 1218 5260 1256
rect 5780 1290 6180 1306
rect 5780 1256 5796 1290
rect 6164 1256 6180 1290
rect 5780 1218 6180 1256
rect 6700 1290 7100 1306
rect 6700 1256 6716 1290
rect 7084 1256 7100 1290
rect 6700 1218 7100 1256
rect 7620 1290 8020 1306
rect 7620 1256 7636 1290
rect 8004 1256 8020 1290
rect 7620 1218 8020 1256
rect 8540 1290 8940 1306
rect 8540 1256 8556 1290
rect 8924 1256 8940 1290
rect 8540 1218 8940 1256
rect -8940 180 -8540 218
rect -8940 146 -8924 180
rect -8556 146 -8540 180
rect -8940 130 -8540 146
rect -8020 180 -7620 218
rect -8020 146 -8004 180
rect -7636 146 -7620 180
rect -8020 130 -7620 146
rect -7100 180 -6700 218
rect -7100 146 -7084 180
rect -6716 146 -6700 180
rect -7100 130 -6700 146
rect -6180 180 -5780 218
rect -6180 146 -6164 180
rect -5796 146 -5780 180
rect -6180 130 -5780 146
rect -5260 180 -4860 218
rect -5260 146 -5244 180
rect -4876 146 -4860 180
rect -5260 130 -4860 146
rect -4340 180 -3940 218
rect -4340 146 -4324 180
rect -3956 146 -3940 180
rect -4340 130 -3940 146
rect -3420 180 -3020 218
rect -3420 146 -3404 180
rect -3036 146 -3020 180
rect -3420 130 -3020 146
rect -2500 180 -2100 218
rect -2500 146 -2484 180
rect -2116 146 -2100 180
rect -2500 130 -2100 146
rect -1580 180 -1180 218
rect -1580 146 -1564 180
rect -1196 146 -1180 180
rect -1580 130 -1180 146
rect -660 180 -260 218
rect -660 146 -644 180
rect -276 146 -260 180
rect -660 130 -260 146
rect 260 180 660 218
rect 260 146 276 180
rect 644 146 660 180
rect 260 130 660 146
rect 1180 180 1580 218
rect 1180 146 1196 180
rect 1564 146 1580 180
rect 1180 130 1580 146
rect 2100 180 2500 218
rect 2100 146 2116 180
rect 2484 146 2500 180
rect 2100 130 2500 146
rect 3020 180 3420 218
rect 3020 146 3036 180
rect 3404 146 3420 180
rect 3020 130 3420 146
rect 3940 180 4340 218
rect 3940 146 3956 180
rect 4324 146 4340 180
rect 3940 130 4340 146
rect 4860 180 5260 218
rect 4860 146 4876 180
rect 5244 146 5260 180
rect 4860 130 5260 146
rect 5780 180 6180 218
rect 5780 146 5796 180
rect 6164 146 6180 180
rect 5780 130 6180 146
rect 6700 180 7100 218
rect 6700 146 6716 180
rect 7084 146 7100 180
rect 6700 130 7100 146
rect 7620 180 8020 218
rect 7620 146 7636 180
rect 8004 146 8020 180
rect 7620 130 8020 146
rect 8540 180 8940 218
rect 8540 146 8556 180
rect 8924 146 8940 180
rect 8540 130 8940 146
rect -8940 -146 -8540 -130
rect -8940 -180 -8924 -146
rect -8556 -180 -8540 -146
rect -8940 -218 -8540 -180
rect -8020 -146 -7620 -130
rect -8020 -180 -8004 -146
rect -7636 -180 -7620 -146
rect -8020 -218 -7620 -180
rect -7100 -146 -6700 -130
rect -7100 -180 -7084 -146
rect -6716 -180 -6700 -146
rect -7100 -218 -6700 -180
rect -6180 -146 -5780 -130
rect -6180 -180 -6164 -146
rect -5796 -180 -5780 -146
rect -6180 -218 -5780 -180
rect -5260 -146 -4860 -130
rect -5260 -180 -5244 -146
rect -4876 -180 -4860 -146
rect -5260 -218 -4860 -180
rect -4340 -146 -3940 -130
rect -4340 -180 -4324 -146
rect -3956 -180 -3940 -146
rect -4340 -218 -3940 -180
rect -3420 -146 -3020 -130
rect -3420 -180 -3404 -146
rect -3036 -180 -3020 -146
rect -3420 -218 -3020 -180
rect -2500 -146 -2100 -130
rect -2500 -180 -2484 -146
rect -2116 -180 -2100 -146
rect -2500 -218 -2100 -180
rect -1580 -146 -1180 -130
rect -1580 -180 -1564 -146
rect -1196 -180 -1180 -146
rect -1580 -218 -1180 -180
rect -660 -146 -260 -130
rect -660 -180 -644 -146
rect -276 -180 -260 -146
rect -660 -218 -260 -180
rect 260 -146 660 -130
rect 260 -180 276 -146
rect 644 -180 660 -146
rect 260 -218 660 -180
rect 1180 -146 1580 -130
rect 1180 -180 1196 -146
rect 1564 -180 1580 -146
rect 1180 -218 1580 -180
rect 2100 -146 2500 -130
rect 2100 -180 2116 -146
rect 2484 -180 2500 -146
rect 2100 -218 2500 -180
rect 3020 -146 3420 -130
rect 3020 -180 3036 -146
rect 3404 -180 3420 -146
rect 3020 -218 3420 -180
rect 3940 -146 4340 -130
rect 3940 -180 3956 -146
rect 4324 -180 4340 -146
rect 3940 -218 4340 -180
rect 4860 -146 5260 -130
rect 4860 -180 4876 -146
rect 5244 -180 5260 -146
rect 4860 -218 5260 -180
rect 5780 -146 6180 -130
rect 5780 -180 5796 -146
rect 6164 -180 6180 -146
rect 5780 -218 6180 -180
rect 6700 -146 7100 -130
rect 6700 -180 6716 -146
rect 7084 -180 7100 -146
rect 6700 -218 7100 -180
rect 7620 -146 8020 -130
rect 7620 -180 7636 -146
rect 8004 -180 8020 -146
rect 7620 -218 8020 -180
rect 8540 -146 8940 -130
rect 8540 -180 8556 -146
rect 8924 -180 8940 -146
rect 8540 -218 8940 -180
rect -8940 -1256 -8540 -1218
rect -8940 -1290 -8924 -1256
rect -8556 -1290 -8540 -1256
rect -8940 -1306 -8540 -1290
rect -8020 -1256 -7620 -1218
rect -8020 -1290 -8004 -1256
rect -7636 -1290 -7620 -1256
rect -8020 -1306 -7620 -1290
rect -7100 -1256 -6700 -1218
rect -7100 -1290 -7084 -1256
rect -6716 -1290 -6700 -1256
rect -7100 -1306 -6700 -1290
rect -6180 -1256 -5780 -1218
rect -6180 -1290 -6164 -1256
rect -5796 -1290 -5780 -1256
rect -6180 -1306 -5780 -1290
rect -5260 -1256 -4860 -1218
rect -5260 -1290 -5244 -1256
rect -4876 -1290 -4860 -1256
rect -5260 -1306 -4860 -1290
rect -4340 -1256 -3940 -1218
rect -4340 -1290 -4324 -1256
rect -3956 -1290 -3940 -1256
rect -4340 -1306 -3940 -1290
rect -3420 -1256 -3020 -1218
rect -3420 -1290 -3404 -1256
rect -3036 -1290 -3020 -1256
rect -3420 -1306 -3020 -1290
rect -2500 -1256 -2100 -1218
rect -2500 -1290 -2484 -1256
rect -2116 -1290 -2100 -1256
rect -2500 -1306 -2100 -1290
rect -1580 -1256 -1180 -1218
rect -1580 -1290 -1564 -1256
rect -1196 -1290 -1180 -1256
rect -1580 -1306 -1180 -1290
rect -660 -1256 -260 -1218
rect -660 -1290 -644 -1256
rect -276 -1290 -260 -1256
rect -660 -1306 -260 -1290
rect 260 -1256 660 -1218
rect 260 -1290 276 -1256
rect 644 -1290 660 -1256
rect 260 -1306 660 -1290
rect 1180 -1256 1580 -1218
rect 1180 -1290 1196 -1256
rect 1564 -1290 1580 -1256
rect 1180 -1306 1580 -1290
rect 2100 -1256 2500 -1218
rect 2100 -1290 2116 -1256
rect 2484 -1290 2500 -1256
rect 2100 -1306 2500 -1290
rect 3020 -1256 3420 -1218
rect 3020 -1290 3036 -1256
rect 3404 -1290 3420 -1256
rect 3020 -1306 3420 -1290
rect 3940 -1256 4340 -1218
rect 3940 -1290 3956 -1256
rect 4324 -1290 4340 -1256
rect 3940 -1306 4340 -1290
rect 4860 -1256 5260 -1218
rect 4860 -1290 4876 -1256
rect 5244 -1290 5260 -1256
rect 4860 -1306 5260 -1290
rect 5780 -1256 6180 -1218
rect 5780 -1290 5796 -1256
rect 6164 -1290 6180 -1256
rect 5780 -1306 6180 -1290
rect 6700 -1256 7100 -1218
rect 6700 -1290 6716 -1256
rect 7084 -1290 7100 -1256
rect 6700 -1306 7100 -1290
rect 7620 -1256 8020 -1218
rect 7620 -1290 7636 -1256
rect 8004 -1290 8020 -1256
rect 7620 -1306 8020 -1290
rect 8540 -1256 8940 -1218
rect 8540 -1290 8556 -1256
rect 8924 -1290 8940 -1256
rect 8540 -1306 8940 -1290
<< polycont >>
rect -8924 1256 -8556 1290
rect -8004 1256 -7636 1290
rect -7084 1256 -6716 1290
rect -6164 1256 -5796 1290
rect -5244 1256 -4876 1290
rect -4324 1256 -3956 1290
rect -3404 1256 -3036 1290
rect -2484 1256 -2116 1290
rect -1564 1256 -1196 1290
rect -644 1256 -276 1290
rect 276 1256 644 1290
rect 1196 1256 1564 1290
rect 2116 1256 2484 1290
rect 3036 1256 3404 1290
rect 3956 1256 4324 1290
rect 4876 1256 5244 1290
rect 5796 1256 6164 1290
rect 6716 1256 7084 1290
rect 7636 1256 8004 1290
rect 8556 1256 8924 1290
rect -8924 146 -8556 180
rect -8004 146 -7636 180
rect -7084 146 -6716 180
rect -6164 146 -5796 180
rect -5244 146 -4876 180
rect -4324 146 -3956 180
rect -3404 146 -3036 180
rect -2484 146 -2116 180
rect -1564 146 -1196 180
rect -644 146 -276 180
rect 276 146 644 180
rect 1196 146 1564 180
rect 2116 146 2484 180
rect 3036 146 3404 180
rect 3956 146 4324 180
rect 4876 146 5244 180
rect 5796 146 6164 180
rect 6716 146 7084 180
rect 7636 146 8004 180
rect 8556 146 8924 180
rect -8924 -180 -8556 -146
rect -8004 -180 -7636 -146
rect -7084 -180 -6716 -146
rect -6164 -180 -5796 -146
rect -5244 -180 -4876 -146
rect -4324 -180 -3956 -146
rect -3404 -180 -3036 -146
rect -2484 -180 -2116 -146
rect -1564 -180 -1196 -146
rect -644 -180 -276 -146
rect 276 -180 644 -146
rect 1196 -180 1564 -146
rect 2116 -180 2484 -146
rect 3036 -180 3404 -146
rect 3956 -180 4324 -146
rect 4876 -180 5244 -146
rect 5796 -180 6164 -146
rect 6716 -180 7084 -146
rect 7636 -180 8004 -146
rect 8556 -180 8924 -146
rect -8924 -1290 -8556 -1256
rect -8004 -1290 -7636 -1256
rect -7084 -1290 -6716 -1256
rect -6164 -1290 -5796 -1256
rect -5244 -1290 -4876 -1256
rect -4324 -1290 -3956 -1256
rect -3404 -1290 -3036 -1256
rect -2484 -1290 -2116 -1256
rect -1564 -1290 -1196 -1256
rect -644 -1290 -276 -1256
rect 276 -1290 644 -1256
rect 1196 -1290 1564 -1256
rect 2116 -1290 2484 -1256
rect 3036 -1290 3404 -1256
rect 3956 -1290 4324 -1256
rect 4876 -1290 5244 -1256
rect 5796 -1290 6164 -1256
rect 6716 -1290 7084 -1256
rect 7636 -1290 8004 -1256
rect 8556 -1290 8924 -1256
<< locali >>
rect -9147 1349 -9051 1383
rect 9051 1349 9147 1383
rect -9147 1287 -9113 1349
rect -8940 1256 -8924 1290
rect -8556 1256 -8540 1290
rect -8020 1256 -8004 1290
rect -7636 1256 -7620 1290
rect -7100 1256 -7084 1290
rect -6716 1256 -6700 1290
rect -6180 1256 -6164 1290
rect -5796 1256 -5780 1290
rect -5260 1256 -5244 1290
rect -4876 1256 -4860 1290
rect -4340 1256 -4324 1290
rect -3956 1256 -3940 1290
rect -3420 1256 -3404 1290
rect -3036 1256 -3020 1290
rect -2500 1256 -2484 1290
rect -2116 1256 -2100 1290
rect -1580 1256 -1564 1290
rect -1196 1256 -1180 1290
rect -660 1256 -644 1290
rect -276 1256 -260 1290
rect 260 1256 276 1290
rect 644 1256 660 1290
rect 1180 1256 1196 1290
rect 1564 1256 1580 1290
rect 2100 1256 2116 1290
rect 2484 1256 2500 1290
rect 3020 1256 3036 1290
rect 3404 1256 3420 1290
rect 3940 1256 3956 1290
rect 4324 1256 4340 1290
rect 4860 1256 4876 1290
rect 5244 1256 5260 1290
rect 5780 1256 5796 1290
rect 6164 1256 6180 1290
rect 6700 1256 6716 1290
rect 7084 1256 7100 1290
rect 7620 1256 7636 1290
rect 8004 1256 8020 1290
rect 8540 1256 8556 1290
rect 8924 1256 8940 1290
rect 9113 1287 9147 1349
rect -9025 1194 -8991 1210
rect -9025 226 -8991 242
rect -8489 1194 -8455 1210
rect -8489 226 -8455 242
rect -8105 1194 -8071 1210
rect -8105 226 -8071 242
rect -7569 1194 -7535 1210
rect -7569 226 -7535 242
rect -7185 1194 -7151 1210
rect -7185 226 -7151 242
rect -6649 1194 -6615 1210
rect -6649 226 -6615 242
rect -6265 1194 -6231 1210
rect -6265 226 -6231 242
rect -5729 1194 -5695 1210
rect -5729 226 -5695 242
rect -5345 1194 -5311 1210
rect -5345 226 -5311 242
rect -4809 1194 -4775 1210
rect -4809 226 -4775 242
rect -4425 1194 -4391 1210
rect -4425 226 -4391 242
rect -3889 1194 -3855 1210
rect -3889 226 -3855 242
rect -3505 1194 -3471 1210
rect -3505 226 -3471 242
rect -2969 1194 -2935 1210
rect -2969 226 -2935 242
rect -2585 1194 -2551 1210
rect -2585 226 -2551 242
rect -2049 1194 -2015 1210
rect -2049 226 -2015 242
rect -1665 1194 -1631 1210
rect -1665 226 -1631 242
rect -1129 1194 -1095 1210
rect -1129 226 -1095 242
rect -745 1194 -711 1210
rect -745 226 -711 242
rect -209 1194 -175 1210
rect -209 226 -175 242
rect 175 1194 209 1210
rect 175 226 209 242
rect 711 1194 745 1210
rect 711 226 745 242
rect 1095 1194 1129 1210
rect 1095 226 1129 242
rect 1631 1194 1665 1210
rect 1631 226 1665 242
rect 2015 1194 2049 1210
rect 2015 226 2049 242
rect 2551 1194 2585 1210
rect 2551 226 2585 242
rect 2935 1194 2969 1210
rect 2935 226 2969 242
rect 3471 1194 3505 1210
rect 3471 226 3505 242
rect 3855 1194 3889 1210
rect 3855 226 3889 242
rect 4391 1194 4425 1210
rect 4391 226 4425 242
rect 4775 1194 4809 1210
rect 4775 226 4809 242
rect 5311 1194 5345 1210
rect 5311 226 5345 242
rect 5695 1194 5729 1210
rect 5695 226 5729 242
rect 6231 1194 6265 1210
rect 6231 226 6265 242
rect 6615 1194 6649 1210
rect 6615 226 6649 242
rect 7151 1194 7185 1210
rect 7151 226 7185 242
rect 7535 1194 7569 1210
rect 7535 226 7569 242
rect 8071 1194 8105 1210
rect 8071 226 8105 242
rect 8455 1194 8489 1210
rect 8455 226 8489 242
rect 8991 1194 9025 1210
rect 8991 226 9025 242
rect -8940 146 -8924 180
rect -8556 146 -8540 180
rect -8020 146 -8004 180
rect -7636 146 -7620 180
rect -7100 146 -7084 180
rect -6716 146 -6700 180
rect -6180 146 -6164 180
rect -5796 146 -5780 180
rect -5260 146 -5244 180
rect -4876 146 -4860 180
rect -4340 146 -4324 180
rect -3956 146 -3940 180
rect -3420 146 -3404 180
rect -3036 146 -3020 180
rect -2500 146 -2484 180
rect -2116 146 -2100 180
rect -1580 146 -1564 180
rect -1196 146 -1180 180
rect -660 146 -644 180
rect -276 146 -260 180
rect 260 146 276 180
rect 644 146 660 180
rect 1180 146 1196 180
rect 1564 146 1580 180
rect 2100 146 2116 180
rect 2484 146 2500 180
rect 3020 146 3036 180
rect 3404 146 3420 180
rect 3940 146 3956 180
rect 4324 146 4340 180
rect 4860 146 4876 180
rect 5244 146 5260 180
rect 5780 146 5796 180
rect 6164 146 6180 180
rect 6700 146 6716 180
rect 7084 146 7100 180
rect 7620 146 7636 180
rect 8004 146 8020 180
rect 8540 146 8556 180
rect 8924 146 8940 180
rect -8940 -180 -8924 -146
rect -8556 -180 -8540 -146
rect -8020 -180 -8004 -146
rect -7636 -180 -7620 -146
rect -7100 -180 -7084 -146
rect -6716 -180 -6700 -146
rect -6180 -180 -6164 -146
rect -5796 -180 -5780 -146
rect -5260 -180 -5244 -146
rect -4876 -180 -4860 -146
rect -4340 -180 -4324 -146
rect -3956 -180 -3940 -146
rect -3420 -180 -3404 -146
rect -3036 -180 -3020 -146
rect -2500 -180 -2484 -146
rect -2116 -180 -2100 -146
rect -1580 -180 -1564 -146
rect -1196 -180 -1180 -146
rect -660 -180 -644 -146
rect -276 -180 -260 -146
rect 260 -180 276 -146
rect 644 -180 660 -146
rect 1180 -180 1196 -146
rect 1564 -180 1580 -146
rect 2100 -180 2116 -146
rect 2484 -180 2500 -146
rect 3020 -180 3036 -146
rect 3404 -180 3420 -146
rect 3940 -180 3956 -146
rect 4324 -180 4340 -146
rect 4860 -180 4876 -146
rect 5244 -180 5260 -146
rect 5780 -180 5796 -146
rect 6164 -180 6180 -146
rect 6700 -180 6716 -146
rect 7084 -180 7100 -146
rect 7620 -180 7636 -146
rect 8004 -180 8020 -146
rect 8540 -180 8556 -146
rect 8924 -180 8940 -146
rect -9025 -242 -8991 -226
rect -9025 -1210 -8991 -1194
rect -8489 -242 -8455 -226
rect -8489 -1210 -8455 -1194
rect -8105 -242 -8071 -226
rect -8105 -1210 -8071 -1194
rect -7569 -242 -7535 -226
rect -7569 -1210 -7535 -1194
rect -7185 -242 -7151 -226
rect -7185 -1210 -7151 -1194
rect -6649 -242 -6615 -226
rect -6649 -1210 -6615 -1194
rect -6265 -242 -6231 -226
rect -6265 -1210 -6231 -1194
rect -5729 -242 -5695 -226
rect -5729 -1210 -5695 -1194
rect -5345 -242 -5311 -226
rect -5345 -1210 -5311 -1194
rect -4809 -242 -4775 -226
rect -4809 -1210 -4775 -1194
rect -4425 -242 -4391 -226
rect -4425 -1210 -4391 -1194
rect -3889 -242 -3855 -226
rect -3889 -1210 -3855 -1194
rect -3505 -242 -3471 -226
rect -3505 -1210 -3471 -1194
rect -2969 -242 -2935 -226
rect -2969 -1210 -2935 -1194
rect -2585 -242 -2551 -226
rect -2585 -1210 -2551 -1194
rect -2049 -242 -2015 -226
rect -2049 -1210 -2015 -1194
rect -1665 -242 -1631 -226
rect -1665 -1210 -1631 -1194
rect -1129 -242 -1095 -226
rect -1129 -1210 -1095 -1194
rect -745 -242 -711 -226
rect -745 -1210 -711 -1194
rect -209 -242 -175 -226
rect -209 -1210 -175 -1194
rect 175 -242 209 -226
rect 175 -1210 209 -1194
rect 711 -242 745 -226
rect 711 -1210 745 -1194
rect 1095 -242 1129 -226
rect 1095 -1210 1129 -1194
rect 1631 -242 1665 -226
rect 1631 -1210 1665 -1194
rect 2015 -242 2049 -226
rect 2015 -1210 2049 -1194
rect 2551 -242 2585 -226
rect 2551 -1210 2585 -1194
rect 2935 -242 2969 -226
rect 2935 -1210 2969 -1194
rect 3471 -242 3505 -226
rect 3471 -1210 3505 -1194
rect 3855 -242 3889 -226
rect 3855 -1210 3889 -1194
rect 4391 -242 4425 -226
rect 4391 -1210 4425 -1194
rect 4775 -242 4809 -226
rect 4775 -1210 4809 -1194
rect 5311 -242 5345 -226
rect 5311 -1210 5345 -1194
rect 5695 -242 5729 -226
rect 5695 -1210 5729 -1194
rect 6231 -242 6265 -226
rect 6231 -1210 6265 -1194
rect 6615 -242 6649 -226
rect 6615 -1210 6649 -1194
rect 7151 -242 7185 -226
rect 7151 -1210 7185 -1194
rect 7535 -242 7569 -226
rect 7535 -1210 7569 -1194
rect 8071 -242 8105 -226
rect 8071 -1210 8105 -1194
rect 8455 -242 8489 -226
rect 8455 -1210 8489 -1194
rect 8991 -242 9025 -226
rect 8991 -1210 9025 -1194
rect -9147 -1349 -9113 -1287
rect -8940 -1290 -8924 -1256
rect -8556 -1290 -8540 -1256
rect -8020 -1290 -8004 -1256
rect -7636 -1290 -7620 -1256
rect -7100 -1290 -7084 -1256
rect -6716 -1290 -6700 -1256
rect -6180 -1290 -6164 -1256
rect -5796 -1290 -5780 -1256
rect -5260 -1290 -5244 -1256
rect -4876 -1290 -4860 -1256
rect -4340 -1290 -4324 -1256
rect -3956 -1290 -3940 -1256
rect -3420 -1290 -3404 -1256
rect -3036 -1290 -3020 -1256
rect -2500 -1290 -2484 -1256
rect -2116 -1290 -2100 -1256
rect -1580 -1290 -1564 -1256
rect -1196 -1290 -1180 -1256
rect -660 -1290 -644 -1256
rect -276 -1290 -260 -1256
rect 260 -1290 276 -1256
rect 644 -1290 660 -1256
rect 1180 -1290 1196 -1256
rect 1564 -1290 1580 -1256
rect 2100 -1290 2116 -1256
rect 2484 -1290 2500 -1256
rect 3020 -1290 3036 -1256
rect 3404 -1290 3420 -1256
rect 3940 -1290 3956 -1256
rect 4324 -1290 4340 -1256
rect 4860 -1290 4876 -1256
rect 5244 -1290 5260 -1256
rect 5780 -1290 5796 -1256
rect 6164 -1290 6180 -1256
rect 6700 -1290 6716 -1256
rect 7084 -1290 7100 -1256
rect 7620 -1290 7636 -1256
rect 8004 -1290 8020 -1256
rect 8540 -1290 8556 -1256
rect 8924 -1290 8940 -1256
rect 9113 -1349 9147 -1287
rect -9147 -1383 -9051 -1349
rect 9051 -1383 9147 -1349
<< viali >>
rect -8924 1256 -8556 1290
rect -8004 1256 -7636 1290
rect -7084 1256 -6716 1290
rect -6164 1256 -5796 1290
rect -5244 1256 -4876 1290
rect -4324 1256 -3956 1290
rect -3404 1256 -3036 1290
rect -2484 1256 -2116 1290
rect -1564 1256 -1196 1290
rect -644 1256 -276 1290
rect 276 1256 644 1290
rect 1196 1256 1564 1290
rect 2116 1256 2484 1290
rect 3036 1256 3404 1290
rect 3956 1256 4324 1290
rect 4876 1256 5244 1290
rect 5796 1256 6164 1290
rect 6716 1256 7084 1290
rect 7636 1256 8004 1290
rect 8556 1256 8924 1290
rect -9025 242 -8991 1194
rect -8489 242 -8455 1194
rect -8105 242 -8071 1194
rect -7569 242 -7535 1194
rect -7185 242 -7151 1194
rect -6649 242 -6615 1194
rect -6265 242 -6231 1194
rect -5729 242 -5695 1194
rect -5345 242 -5311 1194
rect -4809 242 -4775 1194
rect -4425 242 -4391 1194
rect -3889 242 -3855 1194
rect -3505 242 -3471 1194
rect -2969 242 -2935 1194
rect -2585 242 -2551 1194
rect -2049 242 -2015 1194
rect -1665 242 -1631 1194
rect -1129 242 -1095 1194
rect -745 242 -711 1194
rect -209 242 -175 1194
rect 175 242 209 1194
rect 711 242 745 1194
rect 1095 242 1129 1194
rect 1631 242 1665 1194
rect 2015 242 2049 1194
rect 2551 242 2585 1194
rect 2935 242 2969 1194
rect 3471 242 3505 1194
rect 3855 242 3889 1194
rect 4391 242 4425 1194
rect 4775 242 4809 1194
rect 5311 242 5345 1194
rect 5695 242 5729 1194
rect 6231 242 6265 1194
rect 6615 242 6649 1194
rect 7151 242 7185 1194
rect 7535 242 7569 1194
rect 8071 242 8105 1194
rect 8455 242 8489 1194
rect 8991 242 9025 1194
rect -8924 146 -8556 180
rect -8004 146 -7636 180
rect -7084 146 -6716 180
rect -6164 146 -5796 180
rect -5244 146 -4876 180
rect -4324 146 -3956 180
rect -3404 146 -3036 180
rect -2484 146 -2116 180
rect -1564 146 -1196 180
rect -644 146 -276 180
rect 276 146 644 180
rect 1196 146 1564 180
rect 2116 146 2484 180
rect 3036 146 3404 180
rect 3956 146 4324 180
rect 4876 146 5244 180
rect 5796 146 6164 180
rect 6716 146 7084 180
rect 7636 146 8004 180
rect 8556 146 8924 180
rect -8924 -180 -8556 -146
rect -8004 -180 -7636 -146
rect -7084 -180 -6716 -146
rect -6164 -180 -5796 -146
rect -5244 -180 -4876 -146
rect -4324 -180 -3956 -146
rect -3404 -180 -3036 -146
rect -2484 -180 -2116 -146
rect -1564 -180 -1196 -146
rect -644 -180 -276 -146
rect 276 -180 644 -146
rect 1196 -180 1564 -146
rect 2116 -180 2484 -146
rect 3036 -180 3404 -146
rect 3956 -180 4324 -146
rect 4876 -180 5244 -146
rect 5796 -180 6164 -146
rect 6716 -180 7084 -146
rect 7636 -180 8004 -146
rect 8556 -180 8924 -146
rect -9025 -1194 -8991 -242
rect -8489 -1194 -8455 -242
rect -8105 -1194 -8071 -242
rect -7569 -1194 -7535 -242
rect -7185 -1194 -7151 -242
rect -6649 -1194 -6615 -242
rect -6265 -1194 -6231 -242
rect -5729 -1194 -5695 -242
rect -5345 -1194 -5311 -242
rect -4809 -1194 -4775 -242
rect -4425 -1194 -4391 -242
rect -3889 -1194 -3855 -242
rect -3505 -1194 -3471 -242
rect -2969 -1194 -2935 -242
rect -2585 -1194 -2551 -242
rect -2049 -1194 -2015 -242
rect -1665 -1194 -1631 -242
rect -1129 -1194 -1095 -242
rect -745 -1194 -711 -242
rect -209 -1194 -175 -242
rect 175 -1194 209 -242
rect 711 -1194 745 -242
rect 1095 -1194 1129 -242
rect 1631 -1194 1665 -242
rect 2015 -1194 2049 -242
rect 2551 -1194 2585 -242
rect 2935 -1194 2969 -242
rect 3471 -1194 3505 -242
rect 3855 -1194 3889 -242
rect 4391 -1194 4425 -242
rect 4775 -1194 4809 -242
rect 5311 -1194 5345 -242
rect 5695 -1194 5729 -242
rect 6231 -1194 6265 -242
rect 6615 -1194 6649 -242
rect 7151 -1194 7185 -242
rect 7535 -1194 7569 -242
rect 8071 -1194 8105 -242
rect 8455 -1194 8489 -242
rect 8991 -1194 9025 -242
rect -8924 -1290 -8556 -1256
rect -8004 -1290 -7636 -1256
rect -7084 -1290 -6716 -1256
rect -6164 -1290 -5796 -1256
rect -5244 -1290 -4876 -1256
rect -4324 -1290 -3956 -1256
rect -3404 -1290 -3036 -1256
rect -2484 -1290 -2116 -1256
rect -1564 -1290 -1196 -1256
rect -644 -1290 -276 -1256
rect 276 -1290 644 -1256
rect 1196 -1290 1564 -1256
rect 2116 -1290 2484 -1256
rect 3036 -1290 3404 -1256
rect 3956 -1290 4324 -1256
rect 4876 -1290 5244 -1256
rect 5796 -1290 6164 -1256
rect 6716 -1290 7084 -1256
rect 7636 -1290 8004 -1256
rect 8556 -1290 8924 -1256
<< metal1 >>
rect -8936 1290 -8544 1296
rect -8936 1256 -8924 1290
rect -8556 1256 -8544 1290
rect -8936 1250 -8544 1256
rect -8016 1290 -7624 1296
rect -8016 1256 -8004 1290
rect -7636 1256 -7624 1290
rect -8016 1250 -7624 1256
rect -7096 1290 -6704 1296
rect -7096 1256 -7084 1290
rect -6716 1256 -6704 1290
rect -7096 1250 -6704 1256
rect -6176 1290 -5784 1296
rect -6176 1256 -6164 1290
rect -5796 1256 -5784 1290
rect -6176 1250 -5784 1256
rect -5256 1290 -4864 1296
rect -5256 1256 -5244 1290
rect -4876 1256 -4864 1290
rect -5256 1250 -4864 1256
rect -4336 1290 -3944 1296
rect -4336 1256 -4324 1290
rect -3956 1256 -3944 1290
rect -4336 1250 -3944 1256
rect -3416 1290 -3024 1296
rect -3416 1256 -3404 1290
rect -3036 1256 -3024 1290
rect -3416 1250 -3024 1256
rect -2496 1290 -2104 1296
rect -2496 1256 -2484 1290
rect -2116 1256 -2104 1290
rect -2496 1250 -2104 1256
rect -1576 1290 -1184 1296
rect -1576 1256 -1564 1290
rect -1196 1256 -1184 1290
rect -1576 1250 -1184 1256
rect -656 1290 -264 1296
rect -656 1256 -644 1290
rect -276 1256 -264 1290
rect -656 1250 -264 1256
rect 264 1290 656 1296
rect 264 1256 276 1290
rect 644 1256 656 1290
rect 264 1250 656 1256
rect 1184 1290 1576 1296
rect 1184 1256 1196 1290
rect 1564 1256 1576 1290
rect 1184 1250 1576 1256
rect 2104 1290 2496 1296
rect 2104 1256 2116 1290
rect 2484 1256 2496 1290
rect 2104 1250 2496 1256
rect 3024 1290 3416 1296
rect 3024 1256 3036 1290
rect 3404 1256 3416 1290
rect 3024 1250 3416 1256
rect 3944 1290 4336 1296
rect 3944 1256 3956 1290
rect 4324 1256 4336 1290
rect 3944 1250 4336 1256
rect 4864 1290 5256 1296
rect 4864 1256 4876 1290
rect 5244 1256 5256 1290
rect 4864 1250 5256 1256
rect 5784 1290 6176 1296
rect 5784 1256 5796 1290
rect 6164 1256 6176 1290
rect 5784 1250 6176 1256
rect 6704 1290 7096 1296
rect 6704 1256 6716 1290
rect 7084 1256 7096 1290
rect 6704 1250 7096 1256
rect 7624 1290 8016 1296
rect 7624 1256 7636 1290
rect 8004 1256 8016 1290
rect 7624 1250 8016 1256
rect 8544 1290 8936 1296
rect 8544 1256 8556 1290
rect 8924 1256 8936 1290
rect 8544 1250 8936 1256
rect -9031 1194 -8985 1206
rect -9031 242 -9025 1194
rect -8991 242 -8985 1194
rect -9031 230 -8985 242
rect -8495 1194 -8449 1206
rect -8495 242 -8489 1194
rect -8455 242 -8449 1194
rect -8495 230 -8449 242
rect -8111 1194 -8065 1206
rect -8111 242 -8105 1194
rect -8071 242 -8065 1194
rect -8111 230 -8065 242
rect -7575 1194 -7529 1206
rect -7575 242 -7569 1194
rect -7535 242 -7529 1194
rect -7575 230 -7529 242
rect -7191 1194 -7145 1206
rect -7191 242 -7185 1194
rect -7151 242 -7145 1194
rect -7191 230 -7145 242
rect -6655 1194 -6609 1206
rect -6655 242 -6649 1194
rect -6615 242 -6609 1194
rect -6655 230 -6609 242
rect -6271 1194 -6225 1206
rect -6271 242 -6265 1194
rect -6231 242 -6225 1194
rect -6271 230 -6225 242
rect -5735 1194 -5689 1206
rect -5735 242 -5729 1194
rect -5695 242 -5689 1194
rect -5735 230 -5689 242
rect -5351 1194 -5305 1206
rect -5351 242 -5345 1194
rect -5311 242 -5305 1194
rect -5351 230 -5305 242
rect -4815 1194 -4769 1206
rect -4815 242 -4809 1194
rect -4775 242 -4769 1194
rect -4815 230 -4769 242
rect -4431 1194 -4385 1206
rect -4431 242 -4425 1194
rect -4391 242 -4385 1194
rect -4431 230 -4385 242
rect -3895 1194 -3849 1206
rect -3895 242 -3889 1194
rect -3855 242 -3849 1194
rect -3895 230 -3849 242
rect -3511 1194 -3465 1206
rect -3511 242 -3505 1194
rect -3471 242 -3465 1194
rect -3511 230 -3465 242
rect -2975 1194 -2929 1206
rect -2975 242 -2969 1194
rect -2935 242 -2929 1194
rect -2975 230 -2929 242
rect -2591 1194 -2545 1206
rect -2591 242 -2585 1194
rect -2551 242 -2545 1194
rect -2591 230 -2545 242
rect -2055 1194 -2009 1206
rect -2055 242 -2049 1194
rect -2015 242 -2009 1194
rect -2055 230 -2009 242
rect -1671 1194 -1625 1206
rect -1671 242 -1665 1194
rect -1631 242 -1625 1194
rect -1671 230 -1625 242
rect -1135 1194 -1089 1206
rect -1135 242 -1129 1194
rect -1095 242 -1089 1194
rect -1135 230 -1089 242
rect -751 1194 -705 1206
rect -751 242 -745 1194
rect -711 242 -705 1194
rect -751 230 -705 242
rect -215 1194 -169 1206
rect -215 242 -209 1194
rect -175 242 -169 1194
rect -215 230 -169 242
rect 169 1194 215 1206
rect 169 242 175 1194
rect 209 242 215 1194
rect 169 230 215 242
rect 705 1194 751 1206
rect 705 242 711 1194
rect 745 242 751 1194
rect 705 230 751 242
rect 1089 1194 1135 1206
rect 1089 242 1095 1194
rect 1129 242 1135 1194
rect 1089 230 1135 242
rect 1625 1194 1671 1206
rect 1625 242 1631 1194
rect 1665 242 1671 1194
rect 1625 230 1671 242
rect 2009 1194 2055 1206
rect 2009 242 2015 1194
rect 2049 242 2055 1194
rect 2009 230 2055 242
rect 2545 1194 2591 1206
rect 2545 242 2551 1194
rect 2585 242 2591 1194
rect 2545 230 2591 242
rect 2929 1194 2975 1206
rect 2929 242 2935 1194
rect 2969 242 2975 1194
rect 2929 230 2975 242
rect 3465 1194 3511 1206
rect 3465 242 3471 1194
rect 3505 242 3511 1194
rect 3465 230 3511 242
rect 3849 1194 3895 1206
rect 3849 242 3855 1194
rect 3889 242 3895 1194
rect 3849 230 3895 242
rect 4385 1194 4431 1206
rect 4385 242 4391 1194
rect 4425 242 4431 1194
rect 4385 230 4431 242
rect 4769 1194 4815 1206
rect 4769 242 4775 1194
rect 4809 242 4815 1194
rect 4769 230 4815 242
rect 5305 1194 5351 1206
rect 5305 242 5311 1194
rect 5345 242 5351 1194
rect 5305 230 5351 242
rect 5689 1194 5735 1206
rect 5689 242 5695 1194
rect 5729 242 5735 1194
rect 5689 230 5735 242
rect 6225 1194 6271 1206
rect 6225 242 6231 1194
rect 6265 242 6271 1194
rect 6225 230 6271 242
rect 6609 1194 6655 1206
rect 6609 242 6615 1194
rect 6649 242 6655 1194
rect 6609 230 6655 242
rect 7145 1194 7191 1206
rect 7145 242 7151 1194
rect 7185 242 7191 1194
rect 7145 230 7191 242
rect 7529 1194 7575 1206
rect 7529 242 7535 1194
rect 7569 242 7575 1194
rect 7529 230 7575 242
rect 8065 1194 8111 1206
rect 8065 242 8071 1194
rect 8105 242 8111 1194
rect 8065 230 8111 242
rect 8449 1194 8495 1206
rect 8449 242 8455 1194
rect 8489 242 8495 1194
rect 8449 230 8495 242
rect 8985 1194 9031 1206
rect 8985 242 8991 1194
rect 9025 242 9031 1194
rect 8985 230 9031 242
rect -8936 180 -8544 186
rect -8936 146 -8924 180
rect -8556 146 -8544 180
rect -8936 140 -8544 146
rect -8016 180 -7624 186
rect -8016 146 -8004 180
rect -7636 146 -7624 180
rect -8016 140 -7624 146
rect -7096 180 -6704 186
rect -7096 146 -7084 180
rect -6716 146 -6704 180
rect -7096 140 -6704 146
rect -6176 180 -5784 186
rect -6176 146 -6164 180
rect -5796 146 -5784 180
rect -6176 140 -5784 146
rect -5256 180 -4864 186
rect -5256 146 -5244 180
rect -4876 146 -4864 180
rect -5256 140 -4864 146
rect -4336 180 -3944 186
rect -4336 146 -4324 180
rect -3956 146 -3944 180
rect -4336 140 -3944 146
rect -3416 180 -3024 186
rect -3416 146 -3404 180
rect -3036 146 -3024 180
rect -3416 140 -3024 146
rect -2496 180 -2104 186
rect -2496 146 -2484 180
rect -2116 146 -2104 180
rect -2496 140 -2104 146
rect -1576 180 -1184 186
rect -1576 146 -1564 180
rect -1196 146 -1184 180
rect -1576 140 -1184 146
rect -656 180 -264 186
rect -656 146 -644 180
rect -276 146 -264 180
rect -656 140 -264 146
rect 264 180 656 186
rect 264 146 276 180
rect 644 146 656 180
rect 264 140 656 146
rect 1184 180 1576 186
rect 1184 146 1196 180
rect 1564 146 1576 180
rect 1184 140 1576 146
rect 2104 180 2496 186
rect 2104 146 2116 180
rect 2484 146 2496 180
rect 2104 140 2496 146
rect 3024 180 3416 186
rect 3024 146 3036 180
rect 3404 146 3416 180
rect 3024 140 3416 146
rect 3944 180 4336 186
rect 3944 146 3956 180
rect 4324 146 4336 180
rect 3944 140 4336 146
rect 4864 180 5256 186
rect 4864 146 4876 180
rect 5244 146 5256 180
rect 4864 140 5256 146
rect 5784 180 6176 186
rect 5784 146 5796 180
rect 6164 146 6176 180
rect 5784 140 6176 146
rect 6704 180 7096 186
rect 6704 146 6716 180
rect 7084 146 7096 180
rect 6704 140 7096 146
rect 7624 180 8016 186
rect 7624 146 7636 180
rect 8004 146 8016 180
rect 7624 140 8016 146
rect 8544 180 8936 186
rect 8544 146 8556 180
rect 8924 146 8936 180
rect 8544 140 8936 146
rect -8936 -146 -8544 -140
rect -8936 -180 -8924 -146
rect -8556 -180 -8544 -146
rect -8936 -186 -8544 -180
rect -8016 -146 -7624 -140
rect -8016 -180 -8004 -146
rect -7636 -180 -7624 -146
rect -8016 -186 -7624 -180
rect -7096 -146 -6704 -140
rect -7096 -180 -7084 -146
rect -6716 -180 -6704 -146
rect -7096 -186 -6704 -180
rect -6176 -146 -5784 -140
rect -6176 -180 -6164 -146
rect -5796 -180 -5784 -146
rect -6176 -186 -5784 -180
rect -5256 -146 -4864 -140
rect -5256 -180 -5244 -146
rect -4876 -180 -4864 -146
rect -5256 -186 -4864 -180
rect -4336 -146 -3944 -140
rect -4336 -180 -4324 -146
rect -3956 -180 -3944 -146
rect -4336 -186 -3944 -180
rect -3416 -146 -3024 -140
rect -3416 -180 -3404 -146
rect -3036 -180 -3024 -146
rect -3416 -186 -3024 -180
rect -2496 -146 -2104 -140
rect -2496 -180 -2484 -146
rect -2116 -180 -2104 -146
rect -2496 -186 -2104 -180
rect -1576 -146 -1184 -140
rect -1576 -180 -1564 -146
rect -1196 -180 -1184 -146
rect -1576 -186 -1184 -180
rect -656 -146 -264 -140
rect -656 -180 -644 -146
rect -276 -180 -264 -146
rect -656 -186 -264 -180
rect 264 -146 656 -140
rect 264 -180 276 -146
rect 644 -180 656 -146
rect 264 -186 656 -180
rect 1184 -146 1576 -140
rect 1184 -180 1196 -146
rect 1564 -180 1576 -146
rect 1184 -186 1576 -180
rect 2104 -146 2496 -140
rect 2104 -180 2116 -146
rect 2484 -180 2496 -146
rect 2104 -186 2496 -180
rect 3024 -146 3416 -140
rect 3024 -180 3036 -146
rect 3404 -180 3416 -146
rect 3024 -186 3416 -180
rect 3944 -146 4336 -140
rect 3944 -180 3956 -146
rect 4324 -180 4336 -146
rect 3944 -186 4336 -180
rect 4864 -146 5256 -140
rect 4864 -180 4876 -146
rect 5244 -180 5256 -146
rect 4864 -186 5256 -180
rect 5784 -146 6176 -140
rect 5784 -180 5796 -146
rect 6164 -180 6176 -146
rect 5784 -186 6176 -180
rect 6704 -146 7096 -140
rect 6704 -180 6716 -146
rect 7084 -180 7096 -146
rect 6704 -186 7096 -180
rect 7624 -146 8016 -140
rect 7624 -180 7636 -146
rect 8004 -180 8016 -146
rect 7624 -186 8016 -180
rect 8544 -146 8936 -140
rect 8544 -180 8556 -146
rect 8924 -180 8936 -146
rect 8544 -186 8936 -180
rect -9031 -242 -8985 -230
rect -9031 -1194 -9025 -242
rect -8991 -1194 -8985 -242
rect -9031 -1206 -8985 -1194
rect -8495 -242 -8449 -230
rect -8495 -1194 -8489 -242
rect -8455 -1194 -8449 -242
rect -8495 -1206 -8449 -1194
rect -8111 -242 -8065 -230
rect -8111 -1194 -8105 -242
rect -8071 -1194 -8065 -242
rect -8111 -1206 -8065 -1194
rect -7575 -242 -7529 -230
rect -7575 -1194 -7569 -242
rect -7535 -1194 -7529 -242
rect -7575 -1206 -7529 -1194
rect -7191 -242 -7145 -230
rect -7191 -1194 -7185 -242
rect -7151 -1194 -7145 -242
rect -7191 -1206 -7145 -1194
rect -6655 -242 -6609 -230
rect -6655 -1194 -6649 -242
rect -6615 -1194 -6609 -242
rect -6655 -1206 -6609 -1194
rect -6271 -242 -6225 -230
rect -6271 -1194 -6265 -242
rect -6231 -1194 -6225 -242
rect -6271 -1206 -6225 -1194
rect -5735 -242 -5689 -230
rect -5735 -1194 -5729 -242
rect -5695 -1194 -5689 -242
rect -5735 -1206 -5689 -1194
rect -5351 -242 -5305 -230
rect -5351 -1194 -5345 -242
rect -5311 -1194 -5305 -242
rect -5351 -1206 -5305 -1194
rect -4815 -242 -4769 -230
rect -4815 -1194 -4809 -242
rect -4775 -1194 -4769 -242
rect -4815 -1206 -4769 -1194
rect -4431 -242 -4385 -230
rect -4431 -1194 -4425 -242
rect -4391 -1194 -4385 -242
rect -4431 -1206 -4385 -1194
rect -3895 -242 -3849 -230
rect -3895 -1194 -3889 -242
rect -3855 -1194 -3849 -242
rect -3895 -1206 -3849 -1194
rect -3511 -242 -3465 -230
rect -3511 -1194 -3505 -242
rect -3471 -1194 -3465 -242
rect -3511 -1206 -3465 -1194
rect -2975 -242 -2929 -230
rect -2975 -1194 -2969 -242
rect -2935 -1194 -2929 -242
rect -2975 -1206 -2929 -1194
rect -2591 -242 -2545 -230
rect -2591 -1194 -2585 -242
rect -2551 -1194 -2545 -242
rect -2591 -1206 -2545 -1194
rect -2055 -242 -2009 -230
rect -2055 -1194 -2049 -242
rect -2015 -1194 -2009 -242
rect -2055 -1206 -2009 -1194
rect -1671 -242 -1625 -230
rect -1671 -1194 -1665 -242
rect -1631 -1194 -1625 -242
rect -1671 -1206 -1625 -1194
rect -1135 -242 -1089 -230
rect -1135 -1194 -1129 -242
rect -1095 -1194 -1089 -242
rect -1135 -1206 -1089 -1194
rect -751 -242 -705 -230
rect -751 -1194 -745 -242
rect -711 -1194 -705 -242
rect -751 -1206 -705 -1194
rect -215 -242 -169 -230
rect -215 -1194 -209 -242
rect -175 -1194 -169 -242
rect -215 -1206 -169 -1194
rect 169 -242 215 -230
rect 169 -1194 175 -242
rect 209 -1194 215 -242
rect 169 -1206 215 -1194
rect 705 -242 751 -230
rect 705 -1194 711 -242
rect 745 -1194 751 -242
rect 705 -1206 751 -1194
rect 1089 -242 1135 -230
rect 1089 -1194 1095 -242
rect 1129 -1194 1135 -242
rect 1089 -1206 1135 -1194
rect 1625 -242 1671 -230
rect 1625 -1194 1631 -242
rect 1665 -1194 1671 -242
rect 1625 -1206 1671 -1194
rect 2009 -242 2055 -230
rect 2009 -1194 2015 -242
rect 2049 -1194 2055 -242
rect 2009 -1206 2055 -1194
rect 2545 -242 2591 -230
rect 2545 -1194 2551 -242
rect 2585 -1194 2591 -242
rect 2545 -1206 2591 -1194
rect 2929 -242 2975 -230
rect 2929 -1194 2935 -242
rect 2969 -1194 2975 -242
rect 2929 -1206 2975 -1194
rect 3465 -242 3511 -230
rect 3465 -1194 3471 -242
rect 3505 -1194 3511 -242
rect 3465 -1206 3511 -1194
rect 3849 -242 3895 -230
rect 3849 -1194 3855 -242
rect 3889 -1194 3895 -242
rect 3849 -1206 3895 -1194
rect 4385 -242 4431 -230
rect 4385 -1194 4391 -242
rect 4425 -1194 4431 -242
rect 4385 -1206 4431 -1194
rect 4769 -242 4815 -230
rect 4769 -1194 4775 -242
rect 4809 -1194 4815 -242
rect 4769 -1206 4815 -1194
rect 5305 -242 5351 -230
rect 5305 -1194 5311 -242
rect 5345 -1194 5351 -242
rect 5305 -1206 5351 -1194
rect 5689 -242 5735 -230
rect 5689 -1194 5695 -242
rect 5729 -1194 5735 -242
rect 5689 -1206 5735 -1194
rect 6225 -242 6271 -230
rect 6225 -1194 6231 -242
rect 6265 -1194 6271 -242
rect 6225 -1206 6271 -1194
rect 6609 -242 6655 -230
rect 6609 -1194 6615 -242
rect 6649 -1194 6655 -242
rect 6609 -1206 6655 -1194
rect 7145 -242 7191 -230
rect 7145 -1194 7151 -242
rect 7185 -1194 7191 -242
rect 7145 -1206 7191 -1194
rect 7529 -242 7575 -230
rect 7529 -1194 7535 -242
rect 7569 -1194 7575 -242
rect 7529 -1206 7575 -1194
rect 8065 -242 8111 -230
rect 8065 -1194 8071 -242
rect 8105 -1194 8111 -242
rect 8065 -1206 8111 -1194
rect 8449 -242 8495 -230
rect 8449 -1194 8455 -242
rect 8489 -1194 8495 -242
rect 8449 -1206 8495 -1194
rect 8985 -242 9031 -230
rect 8985 -1194 8991 -242
rect 9025 -1194 9031 -242
rect 8985 -1206 9031 -1194
rect -8936 -1256 -8544 -1250
rect -8936 -1290 -8924 -1256
rect -8556 -1290 -8544 -1256
rect -8936 -1296 -8544 -1290
rect -8016 -1256 -7624 -1250
rect -8016 -1290 -8004 -1256
rect -7636 -1290 -7624 -1256
rect -8016 -1296 -7624 -1290
rect -7096 -1256 -6704 -1250
rect -7096 -1290 -7084 -1256
rect -6716 -1290 -6704 -1256
rect -7096 -1296 -6704 -1290
rect -6176 -1256 -5784 -1250
rect -6176 -1290 -6164 -1256
rect -5796 -1290 -5784 -1256
rect -6176 -1296 -5784 -1290
rect -5256 -1256 -4864 -1250
rect -5256 -1290 -5244 -1256
rect -4876 -1290 -4864 -1256
rect -5256 -1296 -4864 -1290
rect -4336 -1256 -3944 -1250
rect -4336 -1290 -4324 -1256
rect -3956 -1290 -3944 -1256
rect -4336 -1296 -3944 -1290
rect -3416 -1256 -3024 -1250
rect -3416 -1290 -3404 -1256
rect -3036 -1290 -3024 -1256
rect -3416 -1296 -3024 -1290
rect -2496 -1256 -2104 -1250
rect -2496 -1290 -2484 -1256
rect -2116 -1290 -2104 -1256
rect -2496 -1296 -2104 -1290
rect -1576 -1256 -1184 -1250
rect -1576 -1290 -1564 -1256
rect -1196 -1290 -1184 -1256
rect -1576 -1296 -1184 -1290
rect -656 -1256 -264 -1250
rect -656 -1290 -644 -1256
rect -276 -1290 -264 -1256
rect -656 -1296 -264 -1290
rect 264 -1256 656 -1250
rect 264 -1290 276 -1256
rect 644 -1290 656 -1256
rect 264 -1296 656 -1290
rect 1184 -1256 1576 -1250
rect 1184 -1290 1196 -1256
rect 1564 -1290 1576 -1256
rect 1184 -1296 1576 -1290
rect 2104 -1256 2496 -1250
rect 2104 -1290 2116 -1256
rect 2484 -1290 2496 -1256
rect 2104 -1296 2496 -1290
rect 3024 -1256 3416 -1250
rect 3024 -1290 3036 -1256
rect 3404 -1290 3416 -1256
rect 3024 -1296 3416 -1290
rect 3944 -1256 4336 -1250
rect 3944 -1290 3956 -1256
rect 4324 -1290 4336 -1256
rect 3944 -1296 4336 -1290
rect 4864 -1256 5256 -1250
rect 4864 -1290 4876 -1256
rect 5244 -1290 5256 -1256
rect 4864 -1296 5256 -1290
rect 5784 -1256 6176 -1250
rect 5784 -1290 5796 -1256
rect 6164 -1290 6176 -1256
rect 5784 -1296 6176 -1290
rect 6704 -1256 7096 -1250
rect 6704 -1290 6716 -1256
rect 7084 -1290 7096 -1256
rect 6704 -1296 7096 -1290
rect 7624 -1256 8016 -1250
rect 7624 -1290 7636 -1256
rect 8004 -1290 8016 -1256
rect 7624 -1296 8016 -1290
rect 8544 -1256 8936 -1250
rect 8544 -1290 8556 -1256
rect 8924 -1290 8936 -1256
rect 8544 -1296 8936 -1290
<< properties >>
string FIXED_BBOX -9130 -1366 9130 1366
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 5 l 2 m 2 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
