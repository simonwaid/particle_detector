magic
tech sky130A
magscale 1 2
timestamp 1647868710
<< pwell >>
rect -325 -719 325 719
<< nmos >>
rect -129 109 -29 509
rect 29 109 129 509
rect -129 -509 -29 -109
rect 29 -509 129 -109
<< ndiff >>
rect -187 497 -129 509
rect -187 121 -175 497
rect -141 121 -129 497
rect -187 109 -129 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 129 497 187 509
rect 129 121 141 497
rect 175 121 187 497
rect 129 109 187 121
rect -187 -121 -129 -109
rect -187 -497 -175 -121
rect -141 -497 -129 -121
rect -187 -509 -129 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 129 -121 187 -109
rect 129 -497 141 -121
rect 175 -497 187 -121
rect 129 -509 187 -497
<< ndiffc >>
rect -175 121 -141 497
rect -17 121 17 497
rect 141 121 175 497
rect -175 -497 -141 -121
rect -17 -497 17 -121
rect 141 -497 175 -121
<< psubdiff >>
rect -289 649 -193 683
rect 193 649 289 683
rect -289 587 -255 649
rect 255 587 289 649
rect -289 -649 -255 -587
rect 255 -649 289 -587
rect -289 -683 -193 -649
rect 193 -683 289 -649
<< psubdiffcont >>
rect -193 649 193 683
rect -289 -587 -255 587
rect 255 -587 289 587
rect -193 -683 193 -649
<< poly >>
rect -129 581 -29 597
rect -129 547 -113 581
rect -45 547 -29 581
rect -129 509 -29 547
rect 29 581 129 597
rect 29 547 45 581
rect 113 547 129 581
rect 29 509 129 547
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect -129 -547 -29 -509
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -509
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 29 -597 129 -581
<< polycont >>
rect -113 547 -45 581
rect 45 547 113 581
rect -113 37 -45 71
rect 45 37 113 71
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect -113 -581 -45 -547
rect 45 -581 113 -547
<< locali >>
rect -289 649 -193 683
rect 193 649 289 683
rect -289 587 -255 649
rect 255 587 289 649
rect -129 547 -113 581
rect -45 547 -29 581
rect 29 547 45 581
rect 113 547 129 581
rect -175 497 -141 513
rect -175 105 -141 121
rect -17 497 17 513
rect -17 105 17 121
rect 141 497 175 513
rect 141 105 175 121
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect -175 -121 -141 -105
rect -175 -513 -141 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 141 -121 175 -105
rect 141 -513 175 -497
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 113 -581 129 -547
rect -289 -649 -255 -587
rect 255 -649 289 -587
rect -289 -683 -193 -649
rect 193 -683 289 -649
<< viali >>
rect -113 547 -45 581
rect 45 547 113 581
rect -175 121 -141 497
rect -17 121 17 497
rect 141 121 175 497
rect -113 37 -45 71
rect 45 37 113 71
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect -175 -497 -141 -121
rect -17 -497 17 -121
rect 141 -497 175 -121
rect -113 -581 -45 -547
rect 45 -581 113 -547
<< metal1 >>
rect -125 581 -33 587
rect -125 547 -113 581
rect -45 547 -33 581
rect -125 541 -33 547
rect 33 581 125 587
rect 33 547 45 581
rect 113 547 125 581
rect 33 541 125 547
rect -181 497 -135 509
rect -181 121 -175 497
rect -141 121 -135 497
rect -181 109 -135 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 135 497 181 509
rect 135 121 141 497
rect 175 121 181 497
rect 135 109 181 121
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect -181 -121 -135 -109
rect -181 -497 -175 -121
rect -141 -497 -135 -121
rect -181 -509 -135 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 135 -121 181 -109
rect 135 -497 141 -121
rect 175 -497 181 -121
rect 135 -509 181 -497
rect -125 -547 -33 -541
rect -125 -581 -113 -547
rect -45 -581 -33 -547
rect -125 -587 -33 -581
rect 33 -547 125 -541
rect 33 -581 45 -547
rect 113 -581 125 -547
rect 33 -587 125 -581
<< properties >>
string FIXED_BBOX -272 -666 272 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.5 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
