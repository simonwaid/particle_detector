magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< poly >>
rect 122 622 476 638
rect 122 588 138 622
rect 172 588 330 622
rect 364 588 476 622
rect 122 572 476 588
rect 122 112 476 128
rect 122 78 234 112
rect 268 78 426 112
rect 460 78 476 112
rect 122 62 476 78
<< polycont >>
rect 138 588 172 622
rect 330 588 364 622
rect 234 78 268 112
rect 426 78 460 112
<< locali >>
rect 122 588 138 622
rect 172 588 330 622
rect 364 588 476 622
rect 122 78 234 112
rect 268 78 426 112
rect 460 78 476 112
rect 80 -100 530 -10
rect 390 -820 500 -100
<< viali >>
rect 138 588 172 622
rect 330 588 364 622
rect 234 78 268 112
rect 426 78 460 112
<< metal1 >>
rect 122 622 476 628
rect 122 620 138 622
rect 0 590 138 620
rect 0 110 30 590
rect 122 588 138 590
rect 172 588 330 622
rect 364 588 476 622
rect 122 582 476 588
rect 164 390 174 550
rect 232 390 242 550
rect 356 390 366 550
rect 424 390 434 550
rect 68 150 78 310
rect 136 150 146 310
rect 260 150 270 310
rect 328 150 338 310
rect 452 150 462 310
rect 520 150 530 310
rect 290 118 320 120
rect 122 112 476 118
rect 122 110 234 112
rect 0 80 234 110
rect 122 78 234 80
rect 268 78 426 112
rect 460 78 476 112
rect 122 72 476 78
rect 130 -420 140 -260
rect 220 -420 230 -260
rect 290 -730 320 72
rect 390 -660 520 -520
rect 420 -830 430 -660
rect 520 -830 530 -660
<< via1 >>
rect 174 390 232 550
rect 366 390 424 550
rect 78 150 136 310
rect 270 150 328 310
rect 462 150 520 310
rect 140 -420 220 -260
rect 430 -830 520 -660
<< metal2 >>
rect 170 550 430 560
rect 170 410 174 550
rect 232 410 366 550
rect 174 380 232 390
rect 424 410 430 550
rect 366 380 424 390
rect 78 310 136 320
rect 270 310 328 320
rect 136 150 270 290
rect 462 310 520 320
rect 328 150 462 290
rect 78 140 520 150
rect 140 -260 220 140
rect 140 -430 220 -420
rect 430 -660 520 -650
rect 430 -840 520 -830
use sky130_fd_pr__nfet_01v8_82JNGJ  sky130_fd_pr__nfet_01v8_82JNGJ_0
timestamp 1654768133
transform 1 0 299 0 1 350
box -359 -410 359 410
use sky130_fd_pr__nfet_01v8_PJG2KG  sky130_fd_pr__nfet_01v8_PJG2KG_0
timestamp 1654768133
transform 1 0 306 0 1 -460
box -246 -410 246 410
<< end >>
