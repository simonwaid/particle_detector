magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< locali >>
rect -8350 40 -8250 3160
rect -7010 40 -6890 3080
rect -5220 40 -5090 3070
rect -3390 40 -3300 3070
rect -2050 2990 -1960 3070
rect -2050 1600 -1660 2990
rect -2050 880 -1960 1600
rect -2050 40 -1820 880
rect 310 10 420 3000
rect 2110 40 2220 3080
rect 3910 40 4020 3080
rect 3720 -1630 3910 -880
rect 4210 -1630 4400 -880
rect 4830 -1630 5110 -890
<< viali >>
rect -9010 -10 -8780 80
rect -7730 -10 -7500 80
rect -2810 -20 -2610 70
<< metal1 >>
rect -6790 3490 -3520 3520
rect -6790 3170 -6300 3490
rect -5830 3170 -4490 3490
rect -4020 3170 -3520 3490
rect -9490 2280 -9410 2720
rect -9180 2590 -8760 3040
rect -8540 2590 -8270 3040
rect -7990 2590 -7980 3040
rect -7830 2600 -7430 3030
rect -7260 2600 -7050 3030
rect -6790 2520 -3520 3170
rect -1540 3480 5630 3520
rect -1540 3160 -910 3480
rect -440 3160 1010 3480
rect 1480 3160 2820 3480
rect 3290 3160 4640 3480
rect 5110 3160 5630 3480
rect -3200 2600 -3190 3030
rect -3050 2600 -3040 3030
rect -2870 2590 -2470 3040
rect -2250 2600 -2240 3030
rect -2150 2600 -2140 3030
rect -1540 2440 5630 3160
rect -8130 2280 -8120 2310
rect -9490 2240 -8120 2280
rect -8130 2230 -8120 2240
rect -8060 2230 -8050 2310
rect -5200 1830 -5190 1850
rect -7060 1500 -6880 1510
rect -7060 1400 -7040 1500
rect -6930 1400 -6880 1500
rect -5240 1470 -5190 1830
rect -5100 1770 -5090 1850
rect -1910 1610 -1900 1710
rect -1810 1680 -1800 1710
rect -1810 1610 -1470 1680
rect -720 1610 -710 1700
rect -560 1690 -550 1700
rect -560 1610 -270 1690
rect -5230 1450 -5190 1470
rect -5160 1430 -5150 1580
rect -5090 1430 -5050 1580
rect -7060 1390 -6880 1400
rect -4250 1290 -4240 1500
rect -4170 1290 -4160 1500
rect -1540 1470 -1470 1610
rect -360 1480 -270 1610
rect 280 1560 290 1640
rect 420 1560 460 1640
rect 410 1440 460 1560
rect 1270 1300 1280 1500
rect 1340 1300 1350 1500
rect 2150 1410 2160 1610
rect 2220 1410 2230 1610
rect 3070 1270 3080 1500
rect 3140 1270 3150 1500
rect 3950 1370 3960 1580
rect 4020 1370 4030 1580
rect 4870 1260 4880 1470
rect 4940 1260 4950 1470
rect -9500 160 -9080 610
rect -8860 160 -8450 610
rect -8150 160 -7740 610
rect -7520 160 -7110 610
rect -3200 150 -2790 610
rect -2560 340 -2150 610
rect -2360 150 -2150 340
rect -9022 80 -8768 86
rect -9030 -10 -9020 80
rect -8780 -10 -8768 80
rect -9022 -16 -8768 -10
rect -7742 80 -7488 86
rect -7742 -10 -7730 80
rect -7500 -10 -7488 80
rect -7742 -16 -7488 -10
rect -2822 70 -2598 76
rect -2822 -20 -2810 70
rect -2610 -20 -2598 70
rect -2822 -26 -2598 -20
rect 1180 -970 1190 -940
rect 1070 -1030 1190 -970
rect 1180 -1040 1190 -1030
rect 1290 -1040 1300 -940
rect 1660 -1090 1670 -960
rect 1750 -1090 1760 -960
<< via1 >>
rect -6300 3170 -5830 3490
rect -4490 3170 -4020 3490
rect -8270 2590 -7990 3040
rect -910 3160 -440 3480
rect 1010 3160 1480 3480
rect 2820 3160 3290 3480
rect 4640 3160 5110 3480
rect -3190 2600 -3050 3030
rect -2240 2600 -2150 3030
rect -8120 2230 -8060 2310
rect -7040 1400 -6930 1500
rect -5190 1770 -5100 1850
rect -1900 1610 -1810 1710
rect -710 1610 -560 1700
rect -5150 1430 -5090 1580
rect -4240 1290 -4170 1500
rect 290 1560 420 1640
rect 1280 1300 1340 1500
rect 2160 1410 2220 1610
rect 3080 1270 3140 1500
rect 3960 1370 4020 1580
rect 4880 1260 4940 1470
rect -9020 -10 -9010 80
rect -9010 -10 -8790 80
rect -7730 -10 -7500 80
rect -2810 -20 -2610 70
rect 1190 -1040 1290 -940
rect 1670 -1090 1750 -960
<< metal2 >>
rect -6300 3490 -5830 3500
rect -6300 3160 -5830 3170
rect -4490 3490 -4020 3500
rect -4490 3160 -4020 3170
rect -910 3480 -440 3490
rect -910 3150 -440 3160
rect 1010 3480 1480 3490
rect 1010 3150 1480 3160
rect 2820 3480 3290 3490
rect 2820 3150 3290 3160
rect 4640 3480 5110 3490
rect 4640 3150 5110 3160
rect -8270 3040 -7990 3050
rect -8270 2580 -7990 2590
rect -3190 3030 -3050 3040
rect -8120 2310 -8060 2320
rect -8120 2220 -8060 2230
rect -4630 2220 -4410 2230
rect -3190 2220 -3050 2600
rect -2240 3030 -2150 3040
rect -1900 2950 -1770 2960
rect -2150 2720 -1900 2950
rect -1900 2710 -1770 2720
rect -2240 2590 -2150 2600
rect -3620 2080 -1810 2220
rect -4630 2070 -4410 2080
rect -5190 1850 -5100 1860
rect -5190 1760 -5100 1770
rect -1900 1710 -1810 2080
rect -6370 1620 -6200 1630
rect -7040 1500 -6930 1510
rect -1900 1600 -1810 1610
rect -710 1820 -600 1830
rect 4570 1720 4710 1730
rect -600 1700 -560 1710
rect -710 1600 -560 1610
rect 290 1640 420 1650
rect -5150 1580 -5090 1590
rect 3900 1630 4020 1640
rect 2160 1610 2220 1620
rect 2100 1600 2160 1610
rect -6370 1450 -6200 1460
rect -5210 1570 -5150 1580
rect -1050 1570 -950 1580
rect -5210 1450 -5150 1460
rect -5150 1420 -5090 1430
rect -4330 1500 -4170 1510
rect -7040 1390 -6930 1400
rect -5620 1390 -5270 1400
rect -1050 1460 -950 1470
rect 1020 1590 1120 1600
rect 1020 1480 1120 1490
rect 1280 1500 1340 1510
rect 290 1450 420 1460
rect 1180 1420 1280 1430
rect 2790 1580 2910 1590
rect 2790 1480 2910 1490
rect 3080 1500 3140 1510
rect 2100 1470 2160 1480
rect -4330 1280 -4170 1290
rect 90 1390 230 1400
rect 1940 1410 2040 1420
rect 2160 1400 2220 1410
rect 1940 1300 2040 1310
rect 2980 1360 3080 1370
rect 4570 1570 4710 1580
rect 3900 1480 3960 1490
rect 4880 1470 4940 1480
rect 1180 1290 1340 1300
rect 90 1280 230 1290
rect -5620 1260 -5270 1270
rect 2980 1260 3140 1270
rect 3720 1360 3840 1370
rect 3960 1360 4020 1370
rect 4820 1410 4880 1420
rect 3720 1260 3840 1270
rect 5210 1420 5350 1430
rect 5210 1270 5350 1280
rect 4820 1260 4880 1270
rect 4880 1250 4940 1260
rect 310 350 640 360
rect -6900 310 310 350
rect -6900 100 -6840 310
rect -9020 80 -8790 90
rect -7730 80 -7500 90
rect -6910 80 -6840 100
rect -9030 -10 -9020 80
rect -8790 -10 -7730 80
rect -7500 -10 -6840 80
rect -9030 -70 -6840 -10
rect -6360 300 -2580 310
rect -6360 -70 -5320 300
rect -9030 -80 -5320 -70
rect -4840 70 -2580 300
rect -4840 -20 -2810 70
rect -2610 -20 -2580 70
rect -4840 -80 -2580 -20
rect -9030 -90 -2580 -80
rect -6910 -100 -2580 -90
rect -2100 40 -270 310
rect 60 40 310 310
rect 640 340 1260 350
rect 1670 340 5740 350
rect 640 310 5740 340
rect 640 40 2020 310
rect 2350 40 3810 310
rect 4140 40 5410 310
rect -2100 30 60 40
rect 310 30 640 40
rect 2020 30 2350 40
rect 3810 30 4140 40
rect 5410 30 5740 40
rect -2100 -100 -40 30
rect 3000 -20 3280 -10
rect -6910 -940 -40 -100
rect 880 -30 1110 -20
rect 880 -240 1110 -230
rect 1360 -30 1590 -20
rect 1360 -240 1590 -230
rect 3000 -270 3280 -260
rect 4910 -30 5190 -20
rect 4910 -280 5190 -270
rect 1190 -340 1290 -330
rect 1190 -940 1290 -460
rect 1660 -530 1750 -520
rect 1660 -960 1750 -650
rect 1660 -1030 1670 -960
rect 1190 -1050 1290 -1040
rect 1670 -1100 1750 -1090
rect 5090 -1630 5520 -1330
rect 2990 -2010 5520 -1630
rect -110 -2020 320 -2010
rect 2790 -2020 5520 -2010
rect 320 -2440 1020 -2140
rect -110 -2470 320 -2460
rect 3220 -2310 5090 -2020
rect 2790 -2470 3220 -2460
rect 5090 -2470 5520 -2460
<< via2 >>
rect -6300 3170 -5830 3490
rect -4490 3170 -4020 3490
rect -910 3160 -440 3480
rect 1010 3160 1480 3480
rect 2820 3160 3290 3480
rect 4640 3160 5110 3480
rect -8270 2590 -7990 3040
rect -8120 2230 -8060 2310
rect -1900 2720 -1770 2950
rect -4630 2080 -4410 2220
rect -5190 1770 -5100 1850
rect -7040 1400 -6930 1500
rect -6370 1460 -6200 1620
rect -710 1700 -600 1820
rect -5210 1460 -5150 1570
rect -5150 1460 -5090 1570
rect -5620 1270 -5270 1390
rect -4330 1290 -4240 1500
rect -4240 1290 -4170 1500
rect -1050 1470 -950 1570
rect 290 1560 420 1580
rect 290 1460 420 1560
rect 1020 1490 1120 1590
rect 2100 1480 2160 1600
rect 2160 1480 2220 1600
rect 2790 1490 2910 1580
rect 3900 1580 4020 1630
rect 90 1290 230 1390
rect 1180 1300 1280 1420
rect 1280 1300 1340 1420
rect 1940 1310 2040 1410
rect 3900 1490 3960 1580
rect 3960 1490 4020 1580
rect 4570 1580 4710 1720
rect 2980 1270 3080 1360
rect 3080 1270 3140 1360
rect 3720 1270 3840 1360
rect 4820 1270 4880 1410
rect 4880 1270 4940 1410
rect 5210 1280 5350 1420
rect -6840 -70 -6360 310
rect -5320 -80 -4840 300
rect -2580 -100 -2100 310
rect -270 40 60 310
rect 310 40 640 350
rect 2020 40 2350 310
rect 3810 40 4140 310
rect 5410 40 5740 310
rect 880 -230 1110 -30
rect 1360 -230 1590 -30
rect 3000 -260 3280 -20
rect 4910 -270 5190 -30
rect 1190 -460 1290 -340
rect 1660 -650 1750 -530
rect -110 -2460 320 -2020
rect 2790 -2460 3220 -2020
rect 5090 -2460 5520 -2020
<< metal3 >>
rect -6310 3490 -5820 3495
rect -6310 3170 -6300 3490
rect -5830 3170 -5820 3490
rect -6310 3165 -5820 3170
rect -4500 3490 -4010 3495
rect -4500 3170 -4490 3490
rect -4020 3170 -4010 3490
rect -4500 3165 -4010 3170
rect -920 3480 -430 3485
rect -920 3160 -910 3480
rect -440 3160 -430 3480
rect -9490 2930 -9300 3160
rect -920 3155 -430 3160
rect 1000 3480 1490 3485
rect 1000 3160 1010 3480
rect 1480 3160 1490 3480
rect 1000 3155 1490 3160
rect 2810 3480 3300 3485
rect 2810 3160 2820 3480
rect 3290 3160 3300 3480
rect 2810 3155 3300 3160
rect 4630 3480 5120 3485
rect 4630 3160 4640 3480
rect 5110 3160 5120 3480
rect 4630 3155 5120 3160
rect -8280 3040 -7980 3045
rect -8280 2590 -8270 3040
rect -7990 2590 -7980 3040
rect -1910 2950 -1760 2955
rect -1910 2720 -1900 2950
rect -1770 2720 -1760 2950
rect -1910 2715 -1760 2720
rect -8280 2585 -7980 2590
rect -1900 2490 -1770 2715
rect -1900 2370 -600 2490
rect -8200 2190 -8190 2360
rect -8070 2315 -8060 2360
rect -8070 2310 -8050 2315
rect -8060 2280 -8050 2310
rect -8060 2230 -6960 2280
rect -8070 2220 -6960 2230
rect -8070 2190 -8060 2220
rect -7030 1505 -6960 2220
rect -4640 2220 -4400 2225
rect -4640 2080 -4630 2220
rect -4410 2080 -2980 2220
rect -4640 2075 -4400 2080
rect -5200 1850 -5090 1855
rect -5200 1770 -5190 1850
rect -5080 1770 -5070 1850
rect -710 1825 -600 2370
rect -720 1820 -590 1825
rect -5200 1765 -5090 1770
rect -720 1700 -710 1820
rect -600 1700 -590 1820
rect -720 1695 -590 1700
rect 4560 1720 4720 1725
rect 3890 1630 4030 1635
rect -6380 1620 -6190 1625
rect -7050 1500 -6920 1505
rect -7050 1400 -7040 1500
rect -6930 1400 -6920 1500
rect -6380 1460 -6370 1620
rect -6200 1570 -6190 1620
rect 2090 1600 2230 1605
rect 1010 1590 1130 1595
rect 280 1580 430 1585
rect -5220 1570 -5080 1575
rect -1060 1570 -940 1575
rect -6200 1490 -5210 1570
rect -6200 1460 -6190 1490
rect -6380 1455 -6190 1460
rect -5220 1460 -5210 1490
rect -5090 1490 -5050 1570
rect -4340 1500 -4160 1505
rect -5090 1460 -5080 1490
rect -5220 1455 -5080 1460
rect -7050 1395 -6920 1400
rect -5630 1390 -5260 1395
rect -4340 1390 -4330 1500
rect -5630 1270 -5620 1390
rect -5270 1310 -4330 1390
rect -5270 1270 -5260 1310
rect -4340 1290 -4330 1310
rect -4170 1390 -4160 1500
rect -1060 1470 -1050 1570
rect -950 1560 -940 1570
rect 280 1560 290 1580
rect -950 1480 290 1560
rect -950 1470 -940 1480
rect -1060 1465 -940 1470
rect 280 1460 290 1480
rect 420 1560 430 1580
rect 420 1480 440 1560
rect 1010 1490 1020 1590
rect 1120 1580 1130 1590
rect 2090 1580 2100 1600
rect 1120 1490 2100 1580
rect 1010 1485 1130 1490
rect 2090 1480 2100 1490
rect 2220 1480 2230 1600
rect 2780 1580 2920 1585
rect 3890 1580 3900 1630
rect 2780 1490 2790 1580
rect 2910 1490 3900 1580
rect 4020 1580 4030 1630
rect 4560 1580 4570 1720
rect 4710 1700 4720 1720
rect 4710 1600 5140 1700
rect 4710 1580 4720 1600
rect 4020 1490 4040 1580
rect 4560 1575 4720 1580
rect 2780 1485 2920 1490
rect 3890 1485 4030 1490
rect 420 1460 430 1480
rect 2090 1475 2230 1480
rect 280 1455 430 1460
rect 1170 1420 1350 1425
rect 80 1390 240 1395
rect -4170 1310 -4140 1390
rect -4170 1290 -4160 1310
rect -4340 1285 -4160 1290
rect 80 1290 90 1390
rect 230 1380 240 1390
rect 1170 1380 1180 1420
rect 230 1300 1180 1380
rect 1340 1380 1350 1420
rect 1930 1410 2050 1415
rect 1340 1300 1360 1380
rect 1930 1310 1940 1410
rect 2040 1360 2050 1410
rect 4810 1410 4950 1415
rect 2970 1360 3150 1365
rect 3710 1360 3850 1365
rect 4810 1360 4820 1410
rect 2040 1310 2980 1360
rect 1930 1305 2980 1310
rect 230 1290 240 1300
rect 1170 1295 1350 1300
rect 80 1285 240 1290
rect 1960 1270 2980 1305
rect 3140 1270 3160 1360
rect 3710 1270 3720 1360
rect 3840 1270 4820 1360
rect 4940 1360 4950 1410
rect 4940 1270 4970 1360
rect -5630 1265 -5260 1270
rect 2970 1265 3150 1270
rect 3710 1265 3850 1270
rect 4810 1265 4950 1270
rect -6900 315 -2240 350
rect -6900 310 -2090 315
rect -6900 100 -6840 310
rect -6910 -70 -6840 100
rect -6360 300 -2580 310
rect -6360 -70 -5320 300
rect -6910 -80 -5320 -70
rect -4840 -80 -2580 300
rect -6910 -100 -2580 -80
rect -2100 100 -2090 310
rect -1990 100 -1820 880
rect 5050 670 5140 1600
rect 1190 570 5140 670
rect 5200 1420 5360 1425
rect 5200 1280 5210 1420
rect 5350 1280 5360 1420
rect 5200 1275 5360 1280
rect 300 350 650 355
rect -280 310 70 315
rect -280 100 -270 310
rect -2100 40 -270 100
rect 60 40 70 310
rect -2100 35 70 40
rect 300 40 310 350
rect 640 40 650 350
rect 300 35 650 40
rect -2100 -100 -40 35
rect -6910 -940 -40 -100
rect 870 -30 1120 -25
rect 870 -230 880 -30
rect 1110 -230 1120 -30
rect 870 -235 1120 -230
rect 1190 -335 1290 570
rect 5200 500 5290 1275
rect 1660 400 5290 500
rect 1350 -30 1600 -25
rect 1350 -230 1360 -30
rect 1590 -230 1600 -30
rect 1350 -235 1600 -230
rect 1180 -340 1300 -335
rect 1180 -460 1190 -340
rect 1290 -460 1300 -340
rect 1180 -465 1300 -460
rect 1660 -525 1760 400
rect 2010 310 2360 315
rect 2010 40 2020 310
rect 2350 40 2360 310
rect 2010 35 2360 40
rect 3800 310 4150 315
rect 3800 40 3810 310
rect 4140 40 4150 310
rect 3800 35 4150 40
rect 5400 310 5750 315
rect 5400 40 5410 310
rect 5740 40 5750 310
rect 5400 35 5750 40
rect 2990 -20 3290 -15
rect 2990 -260 3000 -20
rect 3280 -260 3290 -20
rect 2990 -265 3290 -260
rect 4900 -30 5200 -25
rect 4900 -270 4910 -30
rect 5190 -270 5200 -30
rect 4900 -275 5200 -270
rect 1650 -530 1760 -525
rect 1650 -650 1660 -530
rect 1750 -650 1760 -530
rect 1650 -655 1760 -650
rect -120 -2020 330 -2015
rect -120 -2460 -110 -2020
rect 320 -2460 330 -2020
rect -120 -2465 330 -2460
rect 2780 -2020 3230 -2015
rect 2780 -2460 2790 -2020
rect 3220 -2460 3230 -2020
rect 2780 -2465 3230 -2460
rect 5080 -2020 5530 -2015
rect 5080 -2460 5090 -2020
rect 5520 -2460 5530 -2020
rect 5080 -2465 5530 -2460
<< via3 >>
rect -6300 3170 -5830 3490
rect -4490 3170 -4020 3490
rect -910 3160 -440 3480
rect 1010 3160 1480 3480
rect 2820 3160 3290 3480
rect 4640 3160 5110 3480
rect -8270 2590 -7990 3040
rect -1900 2720 -1770 2950
rect -8190 2310 -8070 2360
rect -8190 2230 -8120 2310
rect -8120 2230 -8070 2310
rect -8190 2190 -8070 2230
rect -5190 1770 -5100 1850
rect -5100 1770 -5080 1850
rect -2580 -100 -2100 310
rect -270 40 60 310
rect 310 40 640 350
rect 880 -230 1110 -30
rect 1360 -230 1590 -30
rect 2020 40 2350 310
rect 3810 40 4140 310
rect 5410 40 5740 310
rect 3000 -260 3280 -20
rect 4910 -270 5190 -30
rect -110 -2460 320 -2020
rect 2790 -2460 3220 -2020
rect 5090 -2460 5520 -2020
<< metal4 >>
rect -6301 3490 -5829 3491
rect -6301 3170 -6300 3490
rect -5830 3170 -5829 3490
rect -6301 3169 -5829 3170
rect -4491 3490 -4019 3491
rect -4491 3170 -4490 3490
rect -4020 3170 -4019 3490
rect -4491 3169 -4019 3170
rect -911 3480 -439 3481
rect -911 3160 -910 3480
rect -440 3160 -439 3480
rect -911 3159 -439 3160
rect 1009 3480 1481 3481
rect 1009 3160 1010 3480
rect 1480 3160 1481 3480
rect 1009 3159 1481 3160
rect 2819 3480 3291 3481
rect 2819 3160 2820 3480
rect 3290 3160 3291 3480
rect 2819 3159 3291 3160
rect 4630 3480 5190 3490
rect 4630 3160 4640 3480
rect 5110 3160 5190 3480
rect -8270 3041 -7590 3050
rect -8271 3040 -7590 3041
rect -8271 2590 -8270 3040
rect -7990 2590 -7590 3040
rect -1901 2950 -1769 2951
rect -2270 2720 -1900 2950
rect -1770 2720 -1769 2950
rect -1901 2719 -1769 2720
rect -8271 2589 -7590 2590
rect -8270 2580 -7590 2589
rect -8191 2360 -8069 2361
rect -8650 2190 -8190 2360
rect -8070 2190 -8069 2360
rect -8191 2189 -8069 2190
rect -7960 1650 -7590 2580
rect -5200 1850 -5070 1860
rect -5200 1770 -5190 1850
rect -5080 1770 -5070 1850
rect -5200 1670 -5070 1770
rect 309 350 641 351
rect -2581 310 -2099 311
rect -2581 -100 -2580 310
rect -2100 -100 -2099 310
rect -271 310 61 311
rect -271 40 -270 310
rect 60 40 61 310
rect -271 39 61 40
rect 309 40 310 350
rect 640 40 641 350
rect 309 39 641 40
rect 2019 40 2020 311
rect 2350 40 2351 311
rect 2019 39 2351 40
rect 3809 40 3810 311
rect 4140 40 4141 311
rect 3809 39 4141 40
rect 2999 -20 3281 -19
rect 1110 -29 1390 -20
rect -2581 -101 -2099 -100
rect 879 -30 1591 -29
rect 879 -230 880 -30
rect 1110 -230 1360 -30
rect 1590 -230 1591 -30
rect 879 -231 1591 -230
rect 1110 -350 1390 -231
rect 2999 -260 3000 -20
rect 3280 -260 3281 -20
rect 2999 -261 3281 -260
rect 4630 -29 5190 3160
rect 5409 40 5410 311
rect 5740 40 5741 311
rect 5409 39 5741 40
rect 4630 -30 5191 -29
rect 3000 -350 3280 -261
rect 4630 -270 4910 -30
rect 5190 -270 5191 -30
rect 4630 -271 5191 -270
rect 4630 -350 5190 -271
rect 4630 -670 4910 -350
rect -111 -2020 321 -2019
rect -111 -2460 -110 -2020
rect 320 -2460 321 -2020
rect -111 -2461 321 -2460
rect 2789 -2020 3221 -2019
rect 2789 -2460 2790 -2020
rect 3220 -2460 3221 -2020
rect 2789 -2461 3221 -2460
rect 5089 -2020 5521 -2019
rect 5089 -2460 5090 -2020
rect 5520 -2460 5521 -2020
rect 5089 -2461 5521 -2460
<< via4 >>
rect -6300 3170 -5830 3490
rect -4490 3170 -4020 3490
rect -910 3160 -440 3480
rect 1010 3160 1480 3480
rect 2820 3160 3290 3480
rect 4640 3160 5110 3480
rect -2580 -100 -2100 310
rect -270 40 60 310
rect 310 40 640 350
rect 2020 310 2350 350
rect 2020 40 2350 310
rect 3810 310 4140 350
rect 3810 40 4140 310
rect 5410 310 5740 350
rect 5410 40 5740 310
rect 1110 -670 1390 -350
rect 3000 -670 3280 -350
rect 4910 -670 5190 -350
rect -110 -2460 320 -2020
rect 2790 -2460 3220 -2020
rect 5090 -2460 5520 -2020
<< metal5 >>
rect -9650 3490 5750 3520
rect -9650 3190 -6300 3490
rect -6324 3170 -6300 3190
rect -5830 3190 -4490 3490
rect -5830 3170 -5806 3190
rect -6324 3146 -5806 3170
rect -4514 3170 -4490 3190
rect -4020 3480 5750 3490
rect -4020 3190 -910 3480
rect -4020 3170 -3996 3190
rect -4514 3146 -3996 3170
rect -934 3160 -910 3190
rect -440 3190 1010 3480
rect -440 3160 -416 3190
rect -934 3136 -416 3160
rect 986 3160 1010 3190
rect 1480 3190 2820 3480
rect 1480 3160 1504 3190
rect 986 3136 1504 3160
rect 2796 3160 2820 3190
rect 3290 3190 4640 3480
rect 3290 3160 3314 3190
rect 2796 3136 3314 3160
rect 4616 3160 4640 3190
rect 5110 3190 5750 3480
rect 5110 3160 5134 3190
rect 4616 3136 5134 3160
rect -3200 350 1260 380
rect -3200 310 310 350
rect -3200 -100 -2580 310
rect -2100 40 -270 310
rect 60 40 310 310
rect 640 340 1260 350
rect 1670 350 5770 380
rect 1670 340 2020 350
rect 640 40 2020 340
rect 2350 40 3810 350
rect 4140 40 5410 350
rect 5740 40 5770 350
rect -2100 20 5770 40
rect -2100 16 664 20
rect 1996 16 2374 20
rect 3786 16 4164 20
rect 5386 16 5764 20
rect -2100 -100 310 16
rect -2604 -124 -2076 -100
rect -210 -1996 310 -100
rect 1086 -330 1414 -326
rect 2976 -330 3304 -326
rect 4886 -330 5214 -326
rect 630 -350 5770 -330
rect 630 -670 1110 -350
rect 1390 -670 3000 -350
rect 3280 -670 4910 -350
rect 5190 -670 5770 -350
rect 630 -690 5770 -670
rect 1086 -694 1414 -690
rect 2976 -694 3304 -690
rect 4886 -694 5214 -690
rect -210 -2020 344 -1996
rect 2766 -2020 3244 -1996
rect 5066 -2020 5544 -1996
rect -210 -2460 -110 -2020
rect 320 -2460 2790 -2020
rect 3220 -2460 5090 -2020
rect 5520 -2460 5770 -2020
rect -134 -2484 344 -2460
rect 2766 -2484 3244 -2460
rect 5066 -2484 5544 -2460
use comp_adv3  comp_adv3_0
timestamp 1654760956
transform 1 0 -5750 0 1 910
box 600 -910 2410 2206
use comp_adv3  comp_adv3_1
timestamp 1654760956
transform 1 0 -7550 0 1 910
box 600 -910 2410 2206
use comp_adv3  comp_adv3_2
timestamp 1654760956
transform 1 0 -240 0 1 910
box 600 -910 2410 2206
use comp_adv3  comp_adv3_3
timestamp 1654760956
transform 1 0 1560 0 1 910
box 600 -910 2410 2206
use comp_adv3  comp_adv3_4
timestamp 1654760956
transform 1 0 3360 0 1 910
box 600 -910 2410 2206
use comp_adv3_di  comp_adv3_di_0
timestamp 1654760956
transform 1 0 -2310 0 1 930
box 300 -930 2682 2106
use comp_to_logic  comp_to_logic_0
timestamp 1654760956
transform 1 0 -570 0 1 -3920
box 890 1440 6340 3910
use sky130_fd_pr__cap_mim_m3_1_H9XL9H  sky130_fd_pr__cap_mim_m3_1_H9XL9H_0
timestamp 1654760956
transform -1 0 -2671 0 -1 2500
box -650 -600 649 600
use sky130_fd_pr__cap_mim_m3_1_H9XL9H  sky130_fd_pr__cap_mim_m3_1_H9XL9H_1
timestamp 1654760956
transform -1 0 -9011 0 -1 2410
box -650 -600 649 600
use sky130_fd_pr__cap_mim_m3_2_MJMGTW  sky130_fd_pr__cap_mim_m3_2_MJMGTW_0
timestamp 1654760956
transform -1 0 -6247 0 -1 -379
box -3351 -2101 3373 2101
use sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL  sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL_0
timestamp 1654760956
transform 1 0 -2672 0 1 1598
box -678 -1598 678 1598
use sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL  sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL_1
timestamp 1654760956
transform 1 0 -8972 0 1 1598
box -678 -1598 678 1598
use sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL  sky130_fd_pr__res_xhigh_po_0p35_Z7KPPL_2
timestamp 1654760956
transform 1 0 -7632 0 1 1598
box -678 -1598 678 1598
<< labels >>
rlabel metal1 -7260 2600 -7050 3030 1 InRef
rlabel metal5 -140 -1730 220 -1310 1 VN
rlabel metal5 -9180 3220 -8810 3470 1 VP
rlabel space 5150 1870 5430 2100 1 OutP
rlabel space 4270 1890 4550 2120 1 OutN
rlabel metal3 -9490 3070 -9300 3160 1 In
rlabel space -4610 1890 -4450 2000 1 Outn_20db
rlabel space -3670 1890 -3560 2010 1 Outp_20db
<< end >>
