magic
tech sky130B
magscale 1 2
timestamp 1654166568
<< locali >>
rect 1450 760 1840 2070
rect 640 750 1840 760
rect 640 670 2640 750
rect 1450 660 2640 670
rect 1450 -40 1530 660
rect 470 -160 2350 -40
rect 470 -170 1970 -160
rect 480 -180 590 -170
rect 480 -320 580 -180
rect 480 -720 590 -320
rect 480 -860 580 -720
rect 480 -870 590 -860
rect 2130 -890 2210 -160
<< metal1 >>
rect 760 1500 2520 1950
rect 740 870 750 1310
rect 1340 870 1350 1310
rect 1930 870 1940 1310
rect 2530 870 2540 1310
rect 540 550 590 560
rect 530 510 590 550
rect 540 500 590 510
rect 1710 500 1770 550
rect 580 -790 650 -250
rect 720 -290 1970 -240
rect 720 -310 760 -290
rect 710 -730 760 -310
rect 720 -750 760 -730
rect 720 -800 1970 -750
<< via1 >>
rect 750 870 1340 1310
rect 1940 870 2530 1310
<< metal2 >>
rect 750 1310 1340 1320
rect 1940 1310 2530 1320
rect 720 870 750 1310
rect 1340 870 1360 1310
rect 510 350 610 520
rect 720 350 1360 870
rect 1900 870 1940 1310
rect 2530 870 2540 1310
rect 1690 350 1790 520
rect 1900 350 2540 870
rect 420 270 710 280
rect 920 180 1340 280
rect 420 100 710 110
rect 820 -50 1340 180
rect 1610 270 1900 280
rect 1610 100 1900 110
rect 1990 -50 2450 280
rect 660 -480 760 -310
rect 820 -490 2450 -50
rect 420 -560 2060 -550
rect 710 -720 1610 -560
rect 1900 -720 2060 -560
rect 420 -730 2060 -720
<< via2 >>
rect 420 110 710 270
rect 1610 110 1900 270
rect 420 -720 710 -560
rect 1610 -720 1900 -560
<< metal3 >>
rect 420 275 710 280
rect 410 270 720 275
rect 410 110 420 270
rect 710 110 720 270
rect 410 105 720 110
rect 1600 270 1910 275
rect 1600 110 1610 270
rect 1900 110 1910 270
rect 1600 105 1910 110
rect 420 -555 710 105
rect 1610 -555 1900 105
rect 410 -560 720 -555
rect 410 -720 420 -560
rect 710 -720 720 -560
rect 410 -725 720 -720
rect 1600 -560 1910 -555
rect 1600 -720 1610 -560
rect 1900 -720 1910 -560
rect 1600 -725 1910 -720
rect 420 -730 710 -725
use currm_comp  currm_comp_0
timestamp 1654072472
transform 1 0 510 0 1 -890
box -80 -40 1670 780
use diffamp_element  diffamp_element_0
timestamp 1654015619
transform 1 0 1060 0 1 -308
box 420 208 1618 1028
use diffamp_element  diffamp_element_1
timestamp 1654015619
transform 1 0 -120 0 1 -308
box 420 208 1618 1028
use sky130_fd_pr__res_xhigh_po_2p85_TY94YJ  sky130_fd_pr__res_xhigh_po_2p85_TY94YJ_0
timestamp 1654072472
transform 1 0 1051 0 1 1408
box -451 -698 451 698
use sky130_fd_pr__res_xhigh_po_2p85_TY94YJ  sky130_fd_pr__res_xhigh_po_2p85_TY94YJ_1
timestamp 1654072472
transform 1 0 2231 0 1 1408
box -451 -698 451 698
<< labels >>
rlabel metal2 510 350 610 520 1 Inp2
rlabel space 1400 240 1450 400 1 Inp
rlabel space 1540 240 1590 400 1 Inn
rlabel metal2 1690 350 1790 520 1 Inn2
rlabel via1 970 1010 1070 1180 1 Outn
rlabel via1 2150 1010 2250 1180 1 Outp
rlabel via2 440 -710 600 -580 1 VN
rlabel metal2 660 -480 760 -310 1 bias
rlabel metal1 1480 1570 1760 1860 1 VP
<< end >>
