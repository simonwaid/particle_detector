magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< pwell >>
rect 748 896 846 906
rect 698 850 846 896
rect 748 840 846 850
rect 890 840 1436 906
rect 710 328 860 396
rect 902 328 1436 396
<< poly >>
rect 748 896 846 906
rect 698 890 846 896
rect 698 856 796 890
rect 830 856 846 890
rect 698 850 846 856
rect 748 840 846 850
rect 890 890 1436 906
rect 890 856 1002 890
rect 1036 856 1194 890
rect 1228 856 1386 890
rect 1420 856 1436 890
rect 890 840 1436 856
rect 710 380 860 396
rect 710 346 726 380
rect 760 346 860 380
rect 710 328 860 346
rect 902 380 1436 396
rect 902 346 918 380
rect 952 346 1098 380
rect 1132 346 1290 380
rect 1324 346 1436 380
rect 902 328 1436 346
<< polycont >>
rect 796 856 830 890
rect 1002 856 1036 890
rect 1194 856 1228 890
rect 1386 856 1420 890
rect 726 346 760 380
rect 918 346 952 380
rect 1098 346 1132 380
rect 1290 346 1324 380
<< locali >>
rect 698 856 796 890
rect 830 856 846 890
rect 890 856 1002 890
rect 1036 856 1194 890
rect 1228 856 1386 890
rect 1420 856 1436 890
rect 470 420 580 830
rect 710 346 726 380
rect 760 346 860 380
rect 902 346 918 380
rect 952 346 1098 380
rect 1132 346 1290 380
rect 1324 346 1436 380
<< viali >>
rect 796 856 830 890
rect 1002 856 1036 890
rect 1194 856 1228 890
rect 1386 856 1420 890
rect 726 346 760 380
rect 918 346 952 380
rect 1098 346 1132 380
rect 1290 346 1324 380
<< metal1 >>
rect 480 896 700 900
rect 480 890 846 896
rect 480 856 796 890
rect 830 856 846 890
rect 480 850 846 856
rect 890 890 1570 900
rect 890 856 1002 890
rect 1036 856 1194 890
rect 1228 856 1386 890
rect 1420 856 1570 890
rect 890 850 1570 856
rect 480 310 520 850
rect 646 660 656 820
rect 710 660 720 820
rect 838 660 848 820
rect 902 660 912 820
rect 1030 660 1040 820
rect 1094 660 1104 820
rect 1222 660 1232 820
rect 1286 660 1296 820
rect 1414 660 1424 820
rect 1478 660 1488 820
rect 550 420 560 580
rect 614 420 624 580
rect 742 420 752 580
rect 806 420 816 580
rect 934 420 944 580
rect 998 420 1008 580
rect 1126 420 1136 580
rect 1190 420 1200 580
rect 1318 420 1328 580
rect 1382 420 1392 580
rect 580 340 620 420
rect 1520 390 1570 850
rect 710 386 750 390
rect 710 380 860 386
rect 710 346 726 380
rect 760 346 860 380
rect 710 340 860 346
rect 900 380 1570 390
rect 900 346 918 380
rect 952 346 1098 380
rect 1132 346 1290 380
rect 1324 346 1570 380
rect 900 340 1570 346
rect 710 310 750 340
rect 480 270 750 310
<< via1 >>
rect 656 660 710 820
rect 848 660 902 820
rect 1040 660 1094 820
rect 1232 660 1286 820
rect 1424 660 1478 820
rect 560 420 614 580
rect 752 420 806 580
rect 944 420 998 580
rect 1136 420 1190 580
rect 1328 420 1382 580
<< metal2 >>
rect 656 820 710 830
rect 656 650 710 660
rect 840 820 1480 830
rect 840 660 848 820
rect 902 660 1040 820
rect 1094 660 1232 820
rect 1286 660 1424 820
rect 1478 660 1480 820
rect 840 650 1480 660
rect 560 580 806 590
rect 614 420 752 580
rect 560 410 806 420
rect 940 580 1382 590
rect 940 420 944 580
rect 998 420 1136 580
rect 1190 420 1328 580
rect 940 410 1382 420
use sky130_fd_pr__nfet_01v8_lvt_DG2JGC  sky130_fd_pr__nfet_01v8_lvt_DG2JGC_0
timestamp 1654768133
transform 1 0 1019 0 1 618
box -599 -410 599 410
<< end >>
