magic
tech sky130A
magscale 1 2
timestamp 1654760956
<< error_p >>
rect -678 272 -620 278
rect -560 272 -502 278
rect -442 272 -384 278
rect -324 272 -266 278
rect -206 272 -148 278
rect -88 272 -30 278
rect 30 272 88 278
rect 148 272 206 278
rect 266 272 324 278
rect 384 272 442 278
rect 502 272 560 278
rect 620 272 678 278
rect -678 238 -666 272
rect -560 238 -548 272
rect -442 238 -430 272
rect -324 238 -312 272
rect -206 238 -194 272
rect -88 238 -76 272
rect 30 238 42 272
rect 148 238 160 272
rect 266 238 278 272
rect 384 238 396 272
rect 502 238 514 272
rect 620 238 632 272
rect -678 232 -620 238
rect -560 232 -502 238
rect -442 232 -384 238
rect -324 232 -266 238
rect -206 232 -148 238
rect -88 232 -30 238
rect 30 232 88 238
rect 148 232 206 238
rect 266 232 324 238
rect 384 232 442 238
rect 502 232 560 238
rect 620 232 678 238
rect -678 -238 -620 -232
rect -560 -238 -502 -232
rect -442 -238 -384 -232
rect -324 -238 -266 -232
rect -206 -238 -148 -232
rect -88 -238 -30 -232
rect 30 -238 88 -232
rect 148 -238 206 -232
rect 266 -238 324 -232
rect 384 -238 442 -232
rect 502 -238 560 -232
rect 620 -238 678 -232
rect -678 -272 -666 -238
rect -560 -272 -548 -238
rect -442 -272 -430 -238
rect -324 -272 -312 -238
rect -206 -272 -194 -238
rect -88 -272 -76 -238
rect 30 -272 42 -238
rect 148 -272 160 -238
rect 266 -272 278 -238
rect 384 -272 396 -238
rect 502 -272 514 -238
rect 620 -272 632 -238
rect -678 -278 -620 -272
rect -560 -278 -502 -272
rect -442 -278 -384 -272
rect -324 -278 -266 -272
rect -206 -278 -148 -272
rect -88 -278 -30 -272
rect 30 -278 88 -272
rect 148 -278 206 -272
rect 266 -278 324 -272
rect 384 -278 442 -272
rect 502 -278 560 -272
rect 620 -278 678 -272
<< pwell >>
rect -875 -410 875 410
<< nmoslvt >>
rect -679 -200 -619 200
rect -561 -200 -501 200
rect -443 -200 -383 200
rect -325 -200 -265 200
rect -207 -200 -147 200
rect -89 -200 -29 200
rect 29 -200 89 200
rect 147 -200 207 200
rect 265 -200 325 200
rect 383 -200 443 200
rect 501 -200 561 200
rect 619 -200 679 200
<< ndiff >>
rect -737 188 -679 200
rect -737 -188 -725 188
rect -691 -188 -679 188
rect -737 -200 -679 -188
rect -619 188 -561 200
rect -619 -188 -607 188
rect -573 -188 -561 188
rect -619 -200 -561 -188
rect -501 188 -443 200
rect -501 -188 -489 188
rect -455 -188 -443 188
rect -501 -200 -443 -188
rect -383 188 -325 200
rect -383 -188 -371 188
rect -337 -188 -325 188
rect -383 -200 -325 -188
rect -265 188 -207 200
rect -265 -188 -253 188
rect -219 -188 -207 188
rect -265 -200 -207 -188
rect -147 188 -89 200
rect -147 -188 -135 188
rect -101 -188 -89 188
rect -147 -200 -89 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 89 188 147 200
rect 89 -188 101 188
rect 135 -188 147 188
rect 89 -200 147 -188
rect 207 188 265 200
rect 207 -188 219 188
rect 253 -188 265 188
rect 207 -200 265 -188
rect 325 188 383 200
rect 325 -188 337 188
rect 371 -188 383 188
rect 325 -200 383 -188
rect 443 188 501 200
rect 443 -188 455 188
rect 489 -188 501 188
rect 443 -200 501 -188
rect 561 188 619 200
rect 561 -188 573 188
rect 607 -188 619 188
rect 561 -200 619 -188
rect 679 188 737 200
rect 679 -188 691 188
rect 725 -188 737 188
rect 679 -200 737 -188
<< ndiffc >>
rect -725 -188 -691 188
rect -607 -188 -573 188
rect -489 -188 -455 188
rect -371 -188 -337 188
rect -253 -188 -219 188
rect -135 -188 -101 188
rect -17 -188 17 188
rect 101 -188 135 188
rect 219 -188 253 188
rect 337 -188 371 188
rect 455 -188 489 188
rect 573 -188 607 188
rect 691 -188 725 188
<< psubdiff >>
rect -839 340 -743 374
rect 743 340 839 374
rect -839 278 -805 340
rect 805 278 839 340
rect -839 -340 -805 -278
rect 805 -340 839 -278
rect -839 -374 -743 -340
rect 743 -374 839 -340
<< psubdiffcont >>
rect -743 340 743 374
rect -839 -278 -805 278
rect 805 -278 839 278
rect -743 -374 743 -340
<< poly >>
rect -682 272 -616 288
rect -682 238 -666 272
rect -632 238 -616 272
rect -682 222 -616 238
rect -564 272 -498 288
rect -564 238 -548 272
rect -514 238 -498 272
rect -564 222 -498 238
rect -446 272 -380 288
rect -446 238 -430 272
rect -396 238 -380 272
rect -446 222 -380 238
rect -328 272 -262 288
rect -328 238 -312 272
rect -278 238 -262 272
rect -328 222 -262 238
rect -210 272 -144 288
rect -210 238 -194 272
rect -160 238 -144 272
rect -210 222 -144 238
rect -92 272 -26 288
rect -92 238 -76 272
rect -42 238 -26 272
rect -92 222 -26 238
rect 26 272 92 288
rect 26 238 42 272
rect 76 238 92 272
rect 26 222 92 238
rect 144 272 210 288
rect 144 238 160 272
rect 194 238 210 272
rect 144 222 210 238
rect 262 272 328 288
rect 262 238 278 272
rect 312 238 328 272
rect 262 222 328 238
rect 380 272 446 288
rect 380 238 396 272
rect 430 238 446 272
rect 380 222 446 238
rect 498 272 564 288
rect 498 238 514 272
rect 548 238 564 272
rect 498 222 564 238
rect 616 272 682 288
rect 616 238 632 272
rect 666 238 682 272
rect 616 222 682 238
rect -679 200 -619 222
rect -561 200 -501 222
rect -443 200 -383 222
rect -325 200 -265 222
rect -207 200 -147 222
rect -89 200 -29 222
rect 29 200 89 222
rect 147 200 207 222
rect 265 200 325 222
rect 383 200 443 222
rect 501 200 561 222
rect 619 200 679 222
rect -679 -222 -619 -200
rect -561 -222 -501 -200
rect -443 -222 -383 -200
rect -325 -222 -265 -200
rect -207 -222 -147 -200
rect -89 -222 -29 -200
rect 29 -222 89 -200
rect 147 -222 207 -200
rect 265 -222 325 -200
rect 383 -222 443 -200
rect 501 -222 561 -200
rect 619 -222 679 -200
rect -682 -238 -616 -222
rect -682 -272 -666 -238
rect -632 -272 -616 -238
rect -682 -288 -616 -272
rect -564 -238 -498 -222
rect -564 -272 -548 -238
rect -514 -272 -498 -238
rect -564 -288 -498 -272
rect -446 -238 -380 -222
rect -446 -272 -430 -238
rect -396 -272 -380 -238
rect -446 -288 -380 -272
rect -328 -238 -262 -222
rect -328 -272 -312 -238
rect -278 -272 -262 -238
rect -328 -288 -262 -272
rect -210 -238 -144 -222
rect -210 -272 -194 -238
rect -160 -272 -144 -238
rect -210 -288 -144 -272
rect -92 -238 -26 -222
rect -92 -272 -76 -238
rect -42 -272 -26 -238
rect -92 -288 -26 -272
rect 26 -238 92 -222
rect 26 -272 42 -238
rect 76 -272 92 -238
rect 26 -288 92 -272
rect 144 -238 210 -222
rect 144 -272 160 -238
rect 194 -272 210 -238
rect 144 -288 210 -272
rect 262 -238 328 -222
rect 262 -272 278 -238
rect 312 -272 328 -238
rect 262 -288 328 -272
rect 380 -238 446 -222
rect 380 -272 396 -238
rect 430 -272 446 -238
rect 380 -288 446 -272
rect 498 -238 564 -222
rect 498 -272 514 -238
rect 548 -272 564 -238
rect 498 -288 564 -272
rect 616 -238 682 -222
rect 616 -272 632 -238
rect 666 -272 682 -238
rect 616 -288 682 -272
<< polycont >>
rect -666 238 -632 272
rect -548 238 -514 272
rect -430 238 -396 272
rect -312 238 -278 272
rect -194 238 -160 272
rect -76 238 -42 272
rect 42 238 76 272
rect 160 238 194 272
rect 278 238 312 272
rect 396 238 430 272
rect 514 238 548 272
rect 632 238 666 272
rect -666 -272 -632 -238
rect -548 -272 -514 -238
rect -430 -272 -396 -238
rect -312 -272 -278 -238
rect -194 -272 -160 -238
rect -76 -272 -42 -238
rect 42 -272 76 -238
rect 160 -272 194 -238
rect 278 -272 312 -238
rect 396 -272 430 -238
rect 514 -272 548 -238
rect 632 -272 666 -238
<< locali >>
rect -839 340 -743 374
rect 743 340 839 374
rect -839 278 -805 340
rect 805 278 839 340
rect -682 238 -666 272
rect -632 238 -616 272
rect -564 238 -548 272
rect -514 238 -498 272
rect -446 238 -430 272
rect -396 238 -380 272
rect -328 238 -312 272
rect -278 238 -262 272
rect -210 238 -194 272
rect -160 238 -144 272
rect -92 238 -76 272
rect -42 238 -26 272
rect 26 238 42 272
rect 76 238 92 272
rect 144 238 160 272
rect 194 238 210 272
rect 262 238 278 272
rect 312 238 328 272
rect 380 238 396 272
rect 430 238 446 272
rect 498 238 514 272
rect 548 238 564 272
rect 616 238 632 272
rect 666 238 682 272
rect -725 188 -691 204
rect -725 -204 -691 -188
rect -607 188 -573 204
rect -607 -204 -573 -188
rect -489 188 -455 204
rect -489 -204 -455 -188
rect -371 188 -337 204
rect -371 -204 -337 -188
rect -253 188 -219 204
rect -253 -204 -219 -188
rect -135 188 -101 204
rect -135 -204 -101 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 101 188 135 204
rect 101 -204 135 -188
rect 219 188 253 204
rect 219 -204 253 -188
rect 337 188 371 204
rect 337 -204 371 -188
rect 455 188 489 204
rect 455 -204 489 -188
rect 573 188 607 204
rect 573 -204 607 -188
rect 691 188 725 204
rect 691 -204 725 -188
rect -682 -272 -666 -238
rect -632 -272 -616 -238
rect -564 -272 -548 -238
rect -514 -272 -498 -238
rect -446 -272 -430 -238
rect -396 -272 -380 -238
rect -328 -272 -312 -238
rect -278 -272 -262 -238
rect -210 -272 -194 -238
rect -160 -272 -144 -238
rect -92 -272 -76 -238
rect -42 -272 -26 -238
rect 26 -272 42 -238
rect 76 -272 92 -238
rect 144 -272 160 -238
rect 194 -272 210 -238
rect 262 -272 278 -238
rect 312 -272 328 -238
rect 380 -272 396 -238
rect 430 -272 446 -238
rect 498 -272 514 -238
rect 548 -272 564 -238
rect 616 -272 632 -238
rect 666 -272 682 -238
rect -839 -340 -805 -278
rect 805 -340 839 -278
rect -839 -374 -743 -340
rect 743 -374 839 -340
<< viali >>
rect -666 238 -632 272
rect -548 238 -514 272
rect -430 238 -396 272
rect -312 238 -278 272
rect -194 238 -160 272
rect -76 238 -42 272
rect 42 238 76 272
rect 160 238 194 272
rect 278 238 312 272
rect 396 238 430 272
rect 514 238 548 272
rect 632 238 666 272
rect -725 -188 -691 188
rect -607 -188 -573 188
rect -489 -188 -455 188
rect -371 -188 -337 188
rect -253 -188 -219 188
rect -135 -188 -101 188
rect -17 -188 17 188
rect 101 -188 135 188
rect 219 -188 253 188
rect 337 -188 371 188
rect 455 -188 489 188
rect 573 -188 607 188
rect 691 -188 725 188
rect -666 -272 -632 -238
rect -548 -272 -514 -238
rect -430 -272 -396 -238
rect -312 -272 -278 -238
rect -194 -272 -160 -238
rect -76 -272 -42 -238
rect 42 -272 76 -238
rect 160 -272 194 -238
rect 278 -272 312 -238
rect 396 -272 430 -238
rect 514 -272 548 -238
rect 632 -272 666 -238
<< metal1 >>
rect -678 272 -620 278
rect -678 238 -666 272
rect -632 238 -620 272
rect -678 232 -620 238
rect -560 272 -502 278
rect -560 238 -548 272
rect -514 238 -502 272
rect -560 232 -502 238
rect -442 272 -384 278
rect -442 238 -430 272
rect -396 238 -384 272
rect -442 232 -384 238
rect -324 272 -266 278
rect -324 238 -312 272
rect -278 238 -266 272
rect -324 232 -266 238
rect -206 272 -148 278
rect -206 238 -194 272
rect -160 238 -148 272
rect -206 232 -148 238
rect -88 272 -30 278
rect -88 238 -76 272
rect -42 238 -30 272
rect -88 232 -30 238
rect 30 272 88 278
rect 30 238 42 272
rect 76 238 88 272
rect 30 232 88 238
rect 148 272 206 278
rect 148 238 160 272
rect 194 238 206 272
rect 148 232 206 238
rect 266 272 324 278
rect 266 238 278 272
rect 312 238 324 272
rect 266 232 324 238
rect 384 272 442 278
rect 384 238 396 272
rect 430 238 442 272
rect 384 232 442 238
rect 502 272 560 278
rect 502 238 514 272
rect 548 238 560 272
rect 502 232 560 238
rect 620 272 678 278
rect 620 238 632 272
rect 666 238 678 272
rect 620 232 678 238
rect -731 188 -685 200
rect -731 -188 -725 188
rect -691 -188 -685 188
rect -731 -200 -685 -188
rect -613 188 -567 200
rect -613 -188 -607 188
rect -573 -188 -567 188
rect -613 -200 -567 -188
rect -495 188 -449 200
rect -495 -188 -489 188
rect -455 -188 -449 188
rect -495 -200 -449 -188
rect -377 188 -331 200
rect -377 -188 -371 188
rect -337 -188 -331 188
rect -377 -200 -331 -188
rect -259 188 -213 200
rect -259 -188 -253 188
rect -219 -188 -213 188
rect -259 -200 -213 -188
rect -141 188 -95 200
rect -141 -188 -135 188
rect -101 -188 -95 188
rect -141 -200 -95 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 95 188 141 200
rect 95 -188 101 188
rect 135 -188 141 188
rect 95 -200 141 -188
rect 213 188 259 200
rect 213 -188 219 188
rect 253 -188 259 188
rect 213 -200 259 -188
rect 331 188 377 200
rect 331 -188 337 188
rect 371 -188 377 188
rect 331 -200 377 -188
rect 449 188 495 200
rect 449 -188 455 188
rect 489 -188 495 188
rect 449 -200 495 -188
rect 567 188 613 200
rect 567 -188 573 188
rect 607 -188 613 188
rect 567 -200 613 -188
rect 685 188 731 200
rect 685 -188 691 188
rect 725 -188 731 188
rect 685 -200 731 -188
rect -678 -238 -620 -232
rect -678 -272 -666 -238
rect -632 -272 -620 -238
rect -678 -278 -620 -272
rect -560 -238 -502 -232
rect -560 -272 -548 -238
rect -514 -272 -502 -238
rect -560 -278 -502 -272
rect -442 -238 -384 -232
rect -442 -272 -430 -238
rect -396 -272 -384 -238
rect -442 -278 -384 -272
rect -324 -238 -266 -232
rect -324 -272 -312 -238
rect -278 -272 -266 -238
rect -324 -278 -266 -272
rect -206 -238 -148 -232
rect -206 -272 -194 -238
rect -160 -272 -148 -238
rect -206 -278 -148 -272
rect -88 -238 -30 -232
rect -88 -272 -76 -238
rect -42 -272 -30 -238
rect -88 -278 -30 -272
rect 30 -238 88 -232
rect 30 -272 42 -238
rect 76 -272 88 -238
rect 30 -278 88 -272
rect 148 -238 206 -232
rect 148 -272 160 -238
rect 194 -272 206 -238
rect 148 -278 206 -272
rect 266 -238 324 -232
rect 266 -272 278 -238
rect 312 -272 324 -238
rect 266 -278 324 -272
rect 384 -238 442 -232
rect 384 -272 396 -238
rect 430 -272 442 -238
rect 384 -278 442 -272
rect 502 -238 560 -232
rect 502 -272 514 -238
rect 548 -272 560 -238
rect 502 -278 560 -272
rect 620 -238 678 -232
rect 620 -272 632 -238
rect 666 -272 678 -238
rect 620 -278 678 -272
<< properties >>
string FIXED_BBOX -822 -357 822 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.3 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
