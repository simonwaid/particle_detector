magic
tech sky130A
magscale 1 2
timestamp 1654768133
<< dnwell >>
rect 5500 1960 7780 3880
<< nwell >>
rect 5420 3674 7860 3960
rect 5420 2166 5706 3674
rect 7574 2166 7860 3674
rect 5420 1880 7860 2166
<< pwell >>
rect 5706 2166 7574 3674
<< nsubdiff >>
rect 5457 3903 7823 3923
rect 5457 3869 5537 3903
rect 7743 3869 7823 3903
rect 5457 3849 7823 3869
rect 5457 3843 5531 3849
rect 5457 1997 5477 3843
rect 5511 1997 5531 3843
rect 7749 3843 7823 3849
rect 5457 1991 5531 1997
rect 7749 1997 7769 3843
rect 7803 1997 7823 3843
rect 7749 1991 7823 1997
rect 5457 1971 7823 1991
rect 5457 1937 5537 1971
rect 7743 1937 7823 1971
rect 5457 1917 7823 1937
<< nsubdiffcont >>
rect 5537 3869 7743 3903
rect 5477 1997 5511 3843
rect 7769 1997 7803 3843
rect 5537 1937 7743 1971
<< poly >>
rect 5923 3500 7361 3516
rect 5923 3466 6037 3500
rect 6071 3466 6233 3500
rect 6267 3466 6429 3500
rect 6463 3466 6625 3500
rect 6659 3466 6821 3500
rect 6855 3466 7017 3500
rect 7051 3466 7213 3500
rect 7247 3466 7361 3500
rect 5923 3450 7361 3466
rect 5923 2990 7361 3006
rect 5923 2956 5939 2990
rect 5973 2956 6135 2990
rect 6169 2956 6331 2990
rect 6365 2956 6527 2990
rect 6561 2956 6723 2990
rect 6757 2956 6919 2990
rect 6953 2956 7115 2990
rect 7149 2956 7311 2990
rect 7345 2956 7361 2990
rect 5923 2940 7361 2956
rect 5923 2882 7361 2898
rect 5923 2848 5939 2882
rect 5973 2848 6135 2882
rect 6169 2848 6331 2882
rect 6365 2848 6527 2882
rect 6561 2848 6723 2882
rect 6757 2848 6919 2882
rect 6953 2848 7115 2882
rect 7149 2848 7311 2882
rect 7345 2848 7361 2882
rect 5923 2832 7361 2848
rect 5923 2372 7361 2388
rect 5923 2338 6037 2372
rect 6071 2338 6233 2372
rect 6267 2338 6429 2372
rect 6463 2338 6625 2372
rect 6659 2338 6821 2372
rect 6855 2338 7017 2372
rect 7051 2338 7213 2372
rect 7247 2338 7361 2372
rect 5923 2322 7361 2338
<< polycont >>
rect 6037 3466 6071 3500
rect 6233 3466 6267 3500
rect 6429 3466 6463 3500
rect 6625 3466 6659 3500
rect 6821 3466 6855 3500
rect 7017 3466 7051 3500
rect 7213 3466 7247 3500
rect 5939 2956 5973 2990
rect 6135 2956 6169 2990
rect 6331 2956 6365 2990
rect 6527 2956 6561 2990
rect 6723 2956 6757 2990
rect 6919 2956 6953 2990
rect 7115 2956 7149 2990
rect 7311 2956 7345 2990
rect 5939 2848 5973 2882
rect 6135 2848 6169 2882
rect 6331 2848 6365 2882
rect 6527 2848 6561 2882
rect 6723 2848 6757 2882
rect 6919 2848 6953 2882
rect 7115 2848 7149 2882
rect 7311 2848 7345 2882
rect 6037 2338 6071 2372
rect 6233 2338 6267 2372
rect 6429 2338 6463 2372
rect 6625 2338 6659 2372
rect 6821 2338 6855 2372
rect 7017 2338 7051 2372
rect 7213 2338 7247 2372
<< locali >>
rect 5477 3869 5537 3903
rect 7743 3869 7803 3903
rect 5477 3843 5511 3869
rect 7769 3843 7803 3869
rect 5923 3466 6037 3500
rect 6071 3466 6233 3500
rect 6267 3466 6429 3500
rect 6463 3466 6625 3500
rect 6659 3466 6821 3500
rect 6855 3466 7017 3500
rect 7051 3466 7213 3500
rect 7247 3466 7361 3500
rect 5923 2956 5939 2990
rect 5973 2956 6135 2990
rect 6169 2956 6331 2990
rect 6365 2956 6527 2990
rect 6561 2956 6723 2990
rect 6757 2956 6919 2990
rect 6953 2956 7115 2990
rect 7149 2956 7311 2990
rect 7345 2956 7361 2990
rect 5923 2848 5939 2882
rect 5973 2848 6135 2882
rect 6169 2848 6331 2882
rect 6365 2848 6527 2882
rect 6561 2848 6723 2882
rect 6757 2848 6919 2882
rect 6953 2848 7115 2882
rect 7149 2848 7311 2882
rect 7345 2848 7361 2882
rect 5923 2338 6037 2372
rect 6071 2338 6233 2372
rect 6267 2338 6429 2372
rect 6463 2338 6625 2372
rect 6659 2338 6821 2372
rect 6855 2338 7017 2372
rect 7051 2338 7213 2372
rect 7247 2338 7361 2372
rect 5477 1971 5511 1997
rect 7769 1971 7803 1997
rect 5477 1937 5537 1971
rect 7743 1937 7803 1971
<< viali >>
rect 6037 3466 6071 3500
rect 6233 3466 6267 3500
rect 6429 3466 6463 3500
rect 6625 3466 6659 3500
rect 6821 3466 6855 3500
rect 7017 3466 7051 3500
rect 7213 3466 7247 3500
rect 5939 2956 5973 2990
rect 6135 2956 6169 2990
rect 6331 2956 6365 2990
rect 6527 2956 6561 2990
rect 6723 2956 6757 2990
rect 6919 2956 6953 2990
rect 7115 2956 7149 2990
rect 7311 2956 7345 2990
rect 5939 2848 5973 2882
rect 6135 2848 6169 2882
rect 6331 2848 6365 2882
rect 6527 2848 6561 2882
rect 6723 2848 6757 2882
rect 6919 2848 6953 2882
rect 7115 2848 7149 2882
rect 7311 2848 7345 2882
rect 6037 2338 6071 2372
rect 6233 2338 6267 2372
rect 6429 2338 6463 2372
rect 6625 2338 6659 2372
rect 6821 2338 6855 2372
rect 7017 2338 7051 2372
rect 7213 2338 7247 2372
<< metal1 >>
rect 5969 4403 5979 4563
rect 6031 4403 6041 4563
rect 6285 4403 6295 4563
rect 6347 4403 6357 4563
rect 6601 4403 6611 4563
rect 6663 4403 6673 4563
rect 6917 4403 6927 4563
rect 6979 4403 6989 4563
rect 7233 4403 7243 4563
rect 7295 4403 7305 4563
rect 5811 4163 5821 4323
rect 5873 4163 5883 4323
rect 6127 4163 6137 4323
rect 6189 4163 6199 4323
rect 6443 4163 6453 4323
rect 6505 4163 6515 4323
rect 6759 4163 6769 4323
rect 6821 4163 6831 4323
rect 7075 4163 7085 4323
rect 7137 4163 7147 4323
rect 7391 4163 7401 4323
rect 7453 4163 7463 4323
rect 5923 3500 7361 3516
rect 5923 3466 6037 3500
rect 6071 3466 6233 3500
rect 6267 3466 6429 3500
rect 6463 3466 6625 3500
rect 6659 3466 6821 3500
rect 6855 3466 7017 3500
rect 7051 3466 7213 3500
rect 7247 3466 7361 3500
rect 5923 3460 7361 3466
rect 5871 3268 5881 3428
rect 5933 3268 5943 3428
rect 6067 3268 6077 3428
rect 6129 3268 6139 3428
rect 6263 3268 6273 3428
rect 6325 3268 6335 3428
rect 6459 3268 6469 3428
rect 6521 3268 6531 3428
rect 6655 3268 6665 3428
rect 6717 3268 6727 3428
rect 6851 3268 6861 3428
rect 6913 3268 6923 3428
rect 7047 3268 7057 3428
rect 7109 3268 7119 3428
rect 7243 3268 7253 3428
rect 7305 3268 7315 3428
rect 5969 3028 5979 3188
rect 6031 3028 6041 3188
rect 6165 3028 6175 3188
rect 6227 3028 6237 3188
rect 6361 3028 6371 3188
rect 6423 3028 6433 3188
rect 6557 3028 6567 3188
rect 6619 3028 6629 3188
rect 6753 3028 6763 3188
rect 6815 3028 6825 3188
rect 6949 3028 6959 3188
rect 7011 3028 7021 3188
rect 7145 3028 7155 3188
rect 7207 3028 7217 3188
rect 7341 3028 7351 3188
rect 7403 3028 7413 3188
rect 5923 2990 7361 2996
rect 5923 2956 5939 2990
rect 5973 2956 6135 2990
rect 6169 2956 6331 2990
rect 6365 2956 6527 2990
rect 6561 2956 6723 2990
rect 6757 2956 6919 2990
rect 6953 2956 7115 2990
rect 7149 2956 7311 2990
rect 7345 2956 7361 2990
rect 5923 2940 7361 2956
rect 5923 2882 7361 2898
rect 5923 2848 5939 2882
rect 5973 2848 6135 2882
rect 6169 2848 6331 2882
rect 6365 2848 6527 2882
rect 6561 2848 6723 2882
rect 6757 2848 6919 2882
rect 6953 2848 7115 2882
rect 7149 2848 7311 2882
rect 7345 2848 7361 2882
rect 5923 2842 7361 2848
rect 5969 2650 5979 2810
rect 6031 2650 6041 2810
rect 6165 2650 6175 2810
rect 6227 2650 6237 2810
rect 6361 2650 6371 2810
rect 6423 2650 6433 2810
rect 6557 2650 6567 2810
rect 6619 2650 6629 2810
rect 6753 2650 6763 2810
rect 6815 2650 6825 2810
rect 6949 2650 6959 2810
rect 7011 2650 7021 2810
rect 7145 2650 7155 2810
rect 7207 2650 7217 2810
rect 7341 2650 7351 2810
rect 7403 2650 7413 2810
rect 5871 2410 5881 2570
rect 5933 2410 5943 2570
rect 6067 2410 6077 2570
rect 6129 2410 6139 2570
rect 6263 2410 6273 2570
rect 6325 2410 6335 2570
rect 6459 2410 6469 2570
rect 6521 2410 6531 2570
rect 6655 2410 6665 2570
rect 6717 2410 6727 2570
rect 6851 2410 6861 2570
rect 6913 2410 6923 2570
rect 7047 2410 7057 2570
rect 7109 2410 7119 2570
rect 7243 2410 7253 2570
rect 7305 2410 7315 2570
rect 5923 2372 7361 2378
rect 5923 2338 6037 2372
rect 6071 2338 6233 2372
rect 6267 2338 6429 2372
rect 6463 2338 6625 2372
rect 6659 2338 6821 2372
rect 6855 2338 7017 2372
rect 7051 2338 7213 2372
rect 7247 2338 7361 2372
rect 5923 2322 7361 2338
<< via1 >>
rect 5979 4403 6031 4563
rect 6295 4403 6347 4563
rect 6611 4403 6663 4563
rect 6927 4403 6979 4563
rect 7243 4403 7295 4563
rect 5821 4163 5873 4323
rect 6137 4163 6189 4323
rect 6453 4163 6505 4323
rect 6769 4163 6821 4323
rect 7085 4163 7137 4323
rect 7401 4163 7453 4323
rect 5881 3268 5933 3428
rect 6077 3268 6129 3428
rect 6273 3268 6325 3428
rect 6469 3268 6521 3428
rect 6665 3268 6717 3428
rect 6861 3268 6913 3428
rect 7057 3268 7109 3428
rect 7253 3268 7305 3428
rect 5979 3028 6031 3188
rect 6175 3028 6227 3188
rect 6371 3028 6423 3188
rect 6567 3028 6619 3188
rect 6763 3028 6815 3188
rect 6959 3028 7011 3188
rect 7155 3028 7207 3188
rect 7351 3028 7403 3188
rect 5979 2650 6031 2810
rect 6175 2650 6227 2810
rect 6371 2650 6423 2810
rect 6567 2650 6619 2810
rect 6763 2650 6815 2810
rect 6959 2650 7011 2810
rect 7155 2650 7207 2810
rect 7351 2650 7403 2810
rect 5881 2410 5933 2570
rect 6077 2410 6129 2570
rect 6273 2410 6325 2570
rect 6469 2410 6521 2570
rect 6665 2410 6717 2570
rect 6861 2410 6913 2570
rect 7057 2410 7109 2570
rect 7253 2410 7305 2570
<< metal2 >>
rect 5979 4563 6031 4573
rect 5979 4393 6031 4403
rect 6295 4563 6347 4573
rect 6295 4393 6347 4403
rect 6611 4563 6663 4573
rect 6611 4393 6663 4403
rect 6927 4563 6979 4573
rect 6927 4393 6979 4403
rect 7243 4563 7295 4573
rect 7243 4393 7295 4403
rect 5821 4323 5873 4333
rect 5821 4153 5873 4163
rect 6137 4323 6189 4333
rect 6137 4153 6189 4163
rect 6453 4323 6505 4333
rect 6453 4153 6505 4163
rect 6769 4323 6821 4333
rect 6769 4153 6821 4163
rect 7085 4323 7137 4333
rect 7085 4153 7137 4163
rect 7401 4323 7453 4333
rect 7401 4153 7453 4163
rect 5881 3428 5933 3438
rect 5881 3258 5933 3268
rect 6077 3428 6129 3438
rect 6077 3258 6129 3268
rect 6273 3428 6325 3438
rect 6273 3258 6325 3268
rect 6469 3428 6521 3438
rect 6469 3258 6521 3268
rect 6665 3428 6717 3438
rect 6665 3258 6717 3268
rect 6861 3428 6913 3438
rect 6861 3258 6913 3268
rect 7057 3428 7109 3438
rect 7057 3258 7109 3268
rect 7253 3428 7305 3438
rect 7253 3258 7305 3268
rect 5979 3188 6031 3198
rect 5979 3018 6031 3028
rect 6175 3188 6227 3198
rect 6175 3018 6227 3028
rect 6371 3188 6423 3198
rect 6371 3018 6423 3028
rect 6567 3188 6619 3198
rect 6567 3018 6619 3028
rect 6763 3188 6815 3198
rect 6763 3018 6815 3028
rect 6959 3188 7011 3198
rect 6959 3018 7011 3028
rect 7155 3188 7207 3198
rect 7155 3018 7207 3028
rect 7351 3188 7403 3198
rect 7351 3018 7403 3028
rect 5979 2810 6031 2820
rect 5979 2640 6031 2650
rect 6175 2810 6227 2820
rect 6175 2640 6227 2650
rect 6371 2810 6423 2820
rect 6371 2640 6423 2650
rect 6567 2810 6619 2820
rect 6567 2640 6619 2650
rect 6763 2810 6815 2820
rect 6763 2640 6815 2650
rect 6959 2810 7011 2820
rect 6959 2640 7011 2650
rect 7155 2810 7207 2820
rect 7155 2640 7207 2650
rect 7351 2810 7403 2820
rect 7351 2640 7403 2650
rect 5881 2570 5933 2580
rect 5881 2400 5933 2410
rect 6077 2570 6129 2580
rect 6077 2400 6129 2410
rect 6273 2570 6325 2580
rect 6273 2400 6325 2410
rect 6469 2570 6521 2580
rect 6469 2400 6521 2410
rect 6665 2570 6717 2580
rect 6665 2400 6717 2410
rect 6861 2570 6913 2580
rect 6861 2400 6913 2410
rect 7057 2570 7109 2580
rect 7057 2400 7109 2410
rect 7253 2570 7305 2580
rect 7253 2400 7305 2410
use sky130_fd_pr__nfet_01v8_lvt_62U3RB  sky130_fd_pr__nfet_01v8_lvt_62U3RB_0
timestamp 1654768133
transform 1 0 6642 0 1 2919
box -902 -719 902 719
use sky130_fd_pr__pfet_01v8_GYVK57  sky130_fd_pr__pfet_01v8_GYVK57_0
timestamp 1654768133
transform 1 0 6637 0 1 4363
box -957 -419 957 419
<< end >>
