magic
tech sky130A
magscale 1 2
timestamp 1645541123
<< metal4 >>
rect -2351 2059 2351 2100
rect -2351 -2059 2095 2059
rect 2331 -2059 2351 2059
rect -2351 -2100 2351 -2059
<< via4 >>
rect 2095 -2059 2331 2059
<< mimcap2 >>
rect -2251 1960 1749 2000
rect -2251 -1960 -2211 1960
rect 1709 -1960 1749 1960
rect -2251 -2000 1749 -1960
<< mimcap2contact >>
rect -2211 -1960 1709 1960
<< metal5 >>
rect 2053 2059 2373 2101
rect -2235 1960 1733 1984
rect -2235 -1960 -2211 1960
rect 1709 -1960 1733 1960
rect -2235 -1984 1733 -1960
rect 2053 -2059 2095 2059
rect 2331 -2059 2373 2059
rect 2053 -2101 2373 -2059
<< properties >>
string FIXED_BBOX -2351 -2100 1849 2100
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
